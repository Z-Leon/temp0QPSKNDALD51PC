library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity	v_message_walign	 is         
port(
   mux_control     : in  std_logic;
	ch_message      : in  std_logic_vector(511 downto 0);
	v_message       : in  std_logic_vector(2047 downto 0);
	v_message_align : out  std_logic_vector(2047 downto 0)
   );	 
end	v_message_walign;
  
architecture rtl of v_message_walign is
   signal ch_message_align :std_logic_vector(2047 downto 0);  
  begin
 ch_message_align(15 downto 0) <= ch_message(3 downto 0) & ch_message(3 downto 0) & ch_message(3 downto 0) & ch_message(3 downto 0);
 ch_message_align(31 downto 16) <= ch_message(7 downto 4) & ch_message(7 downto 4) & ch_message(7 downto 4) & ch_message(7 downto 4);
 ch_message_align(47 downto 32) <= ch_message(11 downto 8) & ch_message(11 downto 8) & ch_message(11 downto 8) & ch_message(11 downto 8);
 ch_message_align(63 downto 48) <= ch_message(15 downto 12) & ch_message(15 downto 12) & ch_message(15 downto 12) & ch_message(15 downto 12);
 ch_message_align(79 downto 64) <= ch_message(19 downto 16) & ch_message(19 downto 16) & ch_message(19 downto 16) & ch_message(19 downto 16);
 ch_message_align(95 downto 80) <= ch_message(23 downto 20) & ch_message(23 downto 20) & ch_message(23 downto 20) & ch_message(23 downto 20);
 ch_message_align(111 downto 96) <= ch_message(27 downto 24) & ch_message(27 downto 24) & ch_message(27 downto 24) & ch_message(27 downto 24);
 ch_message_align(127 downto 112) <= ch_message(31 downto 28) & ch_message(31 downto 28) & ch_message(31 downto 28) & ch_message(31 downto 28);
 ch_message_align(143 downto 128) <= ch_message(35 downto 32) & ch_message(35 downto 32) & ch_message(35 downto 32) & ch_message(35 downto 32);
 ch_message_align(159 downto 144) <= ch_message(39 downto 36) & ch_message(39 downto 36) & ch_message(39 downto 36) & ch_message(39 downto 36);
 ch_message_align(175 downto 160) <= ch_message(43 downto 40) & ch_message(43 downto 40) & ch_message(43 downto 40) & ch_message(43 downto 40);
 ch_message_align(191 downto 176) <= ch_message(47 downto 44) & ch_message(47 downto 44) & ch_message(47 downto 44) & ch_message(47 downto 44);
 ch_message_align(207 downto 192) <= ch_message(51 downto 48) & ch_message(51 downto 48) & ch_message(51 downto 48) & ch_message(51 downto 48);
 ch_message_align(223 downto 208) <= ch_message(55 downto 52) & ch_message(55 downto 52) & ch_message(55 downto 52) & ch_message(55 downto 52);
 ch_message_align(239 downto 224) <= ch_message(59 downto 56) & ch_message(59 downto 56) & ch_message(59 downto 56) & ch_message(59 downto 56);
 ch_message_align(255 downto 240) <= ch_message(63 downto 60) & ch_message(63 downto 60) & ch_message(63 downto 60) & ch_message(63 downto 60);
 ch_message_align(271 downto 256) <= ch_message(67 downto 64) & ch_message(67 downto 64) & ch_message(67 downto 64) & ch_message(67 downto 64);
 ch_message_align(287 downto 272) <= ch_message(71 downto 68) & ch_message(71 downto 68) & ch_message(71 downto 68) & ch_message(71 downto 68);
 ch_message_align(303 downto 288) <= ch_message(75 downto 72) & ch_message(75 downto 72) & ch_message(75 downto 72) & ch_message(75 downto 72);
 ch_message_align(319 downto 304) <= ch_message(79 downto 76) & ch_message(79 downto 76) & ch_message(79 downto 76) & ch_message(79 downto 76);
 ch_message_align(335 downto 320) <= ch_message(83 downto 80) & ch_message(83 downto 80) & ch_message(83 downto 80) & ch_message(83 downto 80);
 ch_message_align(351 downto 336) <= ch_message(87 downto 84) & ch_message(87 downto 84) & ch_message(87 downto 84) & ch_message(87 downto 84);
 ch_message_align(367 downto 352) <= ch_message(91 downto 88) & ch_message(91 downto 88) & ch_message(91 downto 88) & ch_message(91 downto 88);
 ch_message_align(383 downto 368) <= ch_message(95 downto 92) & ch_message(95 downto 92) & ch_message(95 downto 92) & ch_message(95 downto 92);
 ch_message_align(399 downto 384) <= ch_message(99 downto 96) & ch_message(99 downto 96) & ch_message(99 downto 96) & ch_message(99 downto 96);
 ch_message_align(415 downto 400) <= ch_message(103 downto 100) & ch_message(103 downto 100) & ch_message(103 downto 100) & ch_message(103 downto 100);
 ch_message_align(431 downto 416) <= ch_message(107 downto 104) & ch_message(107 downto 104) & ch_message(107 downto 104) & ch_message(107 downto 104);
 ch_message_align(447 downto 432) <= ch_message(111 downto 108) & ch_message(111 downto 108) & ch_message(111 downto 108) & ch_message(111 downto 108);
 ch_message_align(463 downto 448) <= ch_message(115 downto 112) & ch_message(115 downto 112) & ch_message(115 downto 112) & ch_message(115 downto 112);
 ch_message_align(479 downto 464) <= ch_message(119 downto 116) & ch_message(119 downto 116) & ch_message(119 downto 116) & ch_message(119 downto 116);
 ch_message_align(495 downto 480) <= ch_message(123 downto 120) & ch_message(123 downto 120) & ch_message(123 downto 120) & ch_message(123 downto 120);
 ch_message_align(511 downto 496) <= ch_message(127 downto 124) & ch_message(127 downto 124) & ch_message(127 downto 124) & ch_message(127 downto 124);
 ch_message_align(527 downto 512) <= ch_message(131 downto 128) & ch_message(131 downto 128) & ch_message(131 downto 128) & ch_message(131 downto 128);
 ch_message_align(543 downto 528) <= ch_message(135 downto 132) & ch_message(135 downto 132) & ch_message(135 downto 132) & ch_message(135 downto 132);
 ch_message_align(559 downto 544) <= ch_message(139 downto 136) & ch_message(139 downto 136) & ch_message(139 downto 136) & ch_message(139 downto 136);
 ch_message_align(575 downto 560) <= ch_message(143 downto 140) & ch_message(143 downto 140) & ch_message(143 downto 140) & ch_message(143 downto 140);
 ch_message_align(591 downto 576) <= ch_message(147 downto 144) & ch_message(147 downto 144) & ch_message(147 downto 144) & ch_message(147 downto 144);
 ch_message_align(607 downto 592) <= ch_message(151 downto 148) & ch_message(151 downto 148) & ch_message(151 downto 148) & ch_message(151 downto 148);
 ch_message_align(623 downto 608) <= ch_message(155 downto 152) & ch_message(155 downto 152) & ch_message(155 downto 152) & ch_message(155 downto 152);
 ch_message_align(639 downto 624) <= ch_message(159 downto 156) & ch_message(159 downto 156) & ch_message(159 downto 156) & ch_message(159 downto 156);
 ch_message_align(655 downto 640) <= ch_message(163 downto 160) & ch_message(163 downto 160) & ch_message(163 downto 160) & ch_message(163 downto 160);
 ch_message_align(671 downto 656) <= ch_message(167 downto 164) & ch_message(167 downto 164) & ch_message(167 downto 164) & ch_message(167 downto 164);
 ch_message_align(687 downto 672) <= ch_message(171 downto 168) & ch_message(171 downto 168) & ch_message(171 downto 168) & ch_message(171 downto 168);
 ch_message_align(703 downto 688) <= ch_message(175 downto 172) & ch_message(175 downto 172) & ch_message(175 downto 172) & ch_message(175 downto 172);
 ch_message_align(719 downto 704) <= ch_message(179 downto 176) & ch_message(179 downto 176) & ch_message(179 downto 176) & ch_message(179 downto 176);
 ch_message_align(735 downto 720) <= ch_message(183 downto 180) & ch_message(183 downto 180) & ch_message(183 downto 180) & ch_message(183 downto 180);
 ch_message_align(751 downto 736) <= ch_message(187 downto 184) & ch_message(187 downto 184) & ch_message(187 downto 184) & ch_message(187 downto 184);
 ch_message_align(767 downto 752) <= ch_message(191 downto 188) & ch_message(191 downto 188) & ch_message(191 downto 188) & ch_message(191 downto 188);
 ch_message_align(783 downto 768) <= ch_message(195 downto 192) & ch_message(195 downto 192) & ch_message(195 downto 192) & ch_message(195 downto 192);
 ch_message_align(799 downto 784) <= ch_message(199 downto 196) & ch_message(199 downto 196) & ch_message(199 downto 196) & ch_message(199 downto 196);
 ch_message_align(815 downto 800) <= ch_message(203 downto 200) & ch_message(203 downto 200) & ch_message(203 downto 200) & ch_message(203 downto 200);
 ch_message_align(831 downto 816) <= ch_message(207 downto 204) & ch_message(207 downto 204) & ch_message(207 downto 204) & ch_message(207 downto 204);
 ch_message_align(847 downto 832) <= ch_message(211 downto 208) & ch_message(211 downto 208) & ch_message(211 downto 208) & ch_message(211 downto 208);
 ch_message_align(863 downto 848) <= ch_message(215 downto 212) & ch_message(215 downto 212) & ch_message(215 downto 212) & ch_message(215 downto 212);
 ch_message_align(879 downto 864) <= ch_message(219 downto 216) & ch_message(219 downto 216) & ch_message(219 downto 216) & ch_message(219 downto 216);
 ch_message_align(895 downto 880) <= ch_message(223 downto 220) & ch_message(223 downto 220) & ch_message(223 downto 220) & ch_message(223 downto 220);
 ch_message_align(911 downto 896) <= ch_message(227 downto 224) & ch_message(227 downto 224) & ch_message(227 downto 224) & ch_message(227 downto 224);
 ch_message_align(927 downto 912) <= ch_message(231 downto 228) & ch_message(231 downto 228) & ch_message(231 downto 228) & ch_message(231 downto 228);
 ch_message_align(943 downto 928) <= ch_message(235 downto 232) & ch_message(235 downto 232) & ch_message(235 downto 232) & ch_message(235 downto 232);
 ch_message_align(959 downto 944) <= ch_message(239 downto 236) & ch_message(239 downto 236) & ch_message(239 downto 236) & ch_message(239 downto 236);
 ch_message_align(975 downto 960) <= ch_message(243 downto 240) & ch_message(243 downto 240) & ch_message(243 downto 240) & ch_message(243 downto 240);
 ch_message_align(991 downto 976) <= ch_message(247 downto 244) & ch_message(247 downto 244) & ch_message(247 downto 244) & ch_message(247 downto 244);
 ch_message_align(1007 downto 992) <= ch_message(251 downto 248) & ch_message(251 downto 248) & ch_message(251 downto 248) & ch_message(251 downto 248);
 ch_message_align(1023 downto 1008) <= ch_message(255 downto 252) & ch_message(255 downto 252) & ch_message(255 downto 252) & ch_message(255 downto 252);
 ch_message_align(1039 downto 1024) <= ch_message(259 downto 256) & ch_message(259 downto 256) & ch_message(259 downto 256) & ch_message(259 downto 256);
 ch_message_align(1055 downto 1040) <= ch_message(263 downto 260) & ch_message(263 downto 260) & ch_message(263 downto 260) & ch_message(263 downto 260);
 ch_message_align(1071 downto 1056) <= ch_message(267 downto 264) & ch_message(267 downto 264) & ch_message(267 downto 264) & ch_message(267 downto 264);
 ch_message_align(1087 downto 1072) <= ch_message(271 downto 268) & ch_message(271 downto 268) & ch_message(271 downto 268) & ch_message(271 downto 268);
 ch_message_align(1103 downto 1088) <= ch_message(275 downto 272) & ch_message(275 downto 272) & ch_message(275 downto 272) & ch_message(275 downto 272);
 ch_message_align(1119 downto 1104) <= ch_message(279 downto 276) & ch_message(279 downto 276) & ch_message(279 downto 276) & ch_message(279 downto 276);
 ch_message_align(1135 downto 1120) <= ch_message(283 downto 280) & ch_message(283 downto 280) & ch_message(283 downto 280) & ch_message(283 downto 280);
 ch_message_align(1151 downto 1136) <= ch_message(287 downto 284) & ch_message(287 downto 284) & ch_message(287 downto 284) & ch_message(287 downto 284);
 ch_message_align(1167 downto 1152) <= ch_message(291 downto 288) & ch_message(291 downto 288) & ch_message(291 downto 288) & ch_message(291 downto 288);
 ch_message_align(1183 downto 1168) <= ch_message(295 downto 292) & ch_message(295 downto 292) & ch_message(295 downto 292) & ch_message(295 downto 292);
 ch_message_align(1199 downto 1184) <= ch_message(299 downto 296) & ch_message(299 downto 296) & ch_message(299 downto 296) & ch_message(299 downto 296);
 ch_message_align(1215 downto 1200) <= ch_message(303 downto 300) & ch_message(303 downto 300) & ch_message(303 downto 300) & ch_message(303 downto 300);
 ch_message_align(1231 downto 1216) <= ch_message(307 downto 304) & ch_message(307 downto 304) & ch_message(307 downto 304) & ch_message(307 downto 304);
 ch_message_align(1247 downto 1232) <= ch_message(311 downto 308) & ch_message(311 downto 308) & ch_message(311 downto 308) & ch_message(311 downto 308);
 ch_message_align(1263 downto 1248) <= ch_message(315 downto 312) & ch_message(315 downto 312) & ch_message(315 downto 312) & ch_message(315 downto 312);
 ch_message_align(1279 downto 1264) <= ch_message(319 downto 316) & ch_message(319 downto 316) & ch_message(319 downto 316) & ch_message(319 downto 316);
 ch_message_align(1295 downto 1280) <= ch_message(323 downto 320) & ch_message(323 downto 320) & ch_message(323 downto 320) & ch_message(323 downto 320);
 ch_message_align(1311 downto 1296) <= ch_message(327 downto 324) & ch_message(327 downto 324) & ch_message(327 downto 324) & ch_message(327 downto 324);
 ch_message_align(1327 downto 1312) <= ch_message(331 downto 328) & ch_message(331 downto 328) & ch_message(331 downto 328) & ch_message(331 downto 328);
 ch_message_align(1343 downto 1328) <= ch_message(335 downto 332) & ch_message(335 downto 332) & ch_message(335 downto 332) & ch_message(335 downto 332);
 ch_message_align(1359 downto 1344) <= ch_message(339 downto 336) & ch_message(339 downto 336) & ch_message(339 downto 336) & ch_message(339 downto 336);
 ch_message_align(1375 downto 1360) <= ch_message(343 downto 340) & ch_message(343 downto 340) & ch_message(343 downto 340) & ch_message(343 downto 340);
 ch_message_align(1391 downto 1376) <= ch_message(347 downto 344) & ch_message(347 downto 344) & ch_message(347 downto 344) & ch_message(347 downto 344);
 ch_message_align(1407 downto 1392) <= ch_message(351 downto 348) & ch_message(351 downto 348) & ch_message(351 downto 348) & ch_message(351 downto 348);
 ch_message_align(1423 downto 1408) <= ch_message(355 downto 352) & ch_message(355 downto 352) & ch_message(355 downto 352) & ch_message(355 downto 352);
 ch_message_align(1439 downto 1424) <= ch_message(359 downto 356) & ch_message(359 downto 356) & ch_message(359 downto 356) & ch_message(359 downto 356);
 ch_message_align(1455 downto 1440) <= ch_message(363 downto 360) & ch_message(363 downto 360) & ch_message(363 downto 360) & ch_message(363 downto 360);
 ch_message_align(1471 downto 1456) <= ch_message(367 downto 364) & ch_message(367 downto 364) & ch_message(367 downto 364) & ch_message(367 downto 364);
 ch_message_align(1487 downto 1472) <= ch_message(371 downto 368) & ch_message(371 downto 368) & ch_message(371 downto 368) & ch_message(371 downto 368);
 ch_message_align(1503 downto 1488) <= ch_message(375 downto 372) & ch_message(375 downto 372) & ch_message(375 downto 372) & ch_message(375 downto 372);
 ch_message_align(1519 downto 1504) <= ch_message(379 downto 376) & ch_message(379 downto 376) & ch_message(379 downto 376) & ch_message(379 downto 376);
 ch_message_align(1535 downto 1520) <= ch_message(383 downto 380) & ch_message(383 downto 380) & ch_message(383 downto 380) & ch_message(383 downto 380);
 ch_message_align(1551 downto 1536) <= ch_message(387 downto 384) & ch_message(387 downto 384) & ch_message(387 downto 384) & ch_message(387 downto 384);
 ch_message_align(1567 downto 1552) <= ch_message(391 downto 388) & ch_message(391 downto 388) & ch_message(391 downto 388) & ch_message(391 downto 388);
 ch_message_align(1583 downto 1568) <= ch_message(395 downto 392) & ch_message(395 downto 392) & ch_message(395 downto 392) & ch_message(395 downto 392);
 ch_message_align(1599 downto 1584) <= ch_message(399 downto 396) & ch_message(399 downto 396) & ch_message(399 downto 396) & ch_message(399 downto 396);
 ch_message_align(1615 downto 1600) <= ch_message(403 downto 400) & ch_message(403 downto 400) & ch_message(403 downto 400) & ch_message(403 downto 400);
 ch_message_align(1631 downto 1616) <= ch_message(407 downto 404) & ch_message(407 downto 404) & ch_message(407 downto 404) & ch_message(407 downto 404);
 ch_message_align(1647 downto 1632) <= ch_message(411 downto 408) & ch_message(411 downto 408) & ch_message(411 downto 408) & ch_message(411 downto 408);
 ch_message_align(1663 downto 1648) <= ch_message(415 downto 412) & ch_message(415 downto 412) & ch_message(415 downto 412) & ch_message(415 downto 412);
 ch_message_align(1679 downto 1664) <= ch_message(419 downto 416) & ch_message(419 downto 416) & ch_message(419 downto 416) & ch_message(419 downto 416);
 ch_message_align(1695 downto 1680) <= ch_message(423 downto 420) & ch_message(423 downto 420) & ch_message(423 downto 420) & ch_message(423 downto 420);
 ch_message_align(1711 downto 1696) <= ch_message(427 downto 424) & ch_message(427 downto 424) & ch_message(427 downto 424) & ch_message(427 downto 424);
 ch_message_align(1727 downto 1712) <= ch_message(431 downto 428) & ch_message(431 downto 428) & ch_message(431 downto 428) & ch_message(431 downto 428);
 ch_message_align(1743 downto 1728) <= ch_message(435 downto 432) & ch_message(435 downto 432) & ch_message(435 downto 432) & ch_message(435 downto 432);
 ch_message_align(1759 downto 1744) <= ch_message(439 downto 436) & ch_message(439 downto 436) & ch_message(439 downto 436) & ch_message(439 downto 436);
 ch_message_align(1775 downto 1760) <= ch_message(443 downto 440) & ch_message(443 downto 440) & ch_message(443 downto 440) & ch_message(443 downto 440);
 ch_message_align(1791 downto 1776) <= ch_message(447 downto 444) & ch_message(447 downto 444) & ch_message(447 downto 444) & ch_message(447 downto 444);
 ch_message_align(1807 downto 1792) <= ch_message(451 downto 448) & ch_message(451 downto 448) & ch_message(451 downto 448) & ch_message(451 downto 448);
 ch_message_align(1823 downto 1808) <= ch_message(455 downto 452) & ch_message(455 downto 452) & ch_message(455 downto 452) & ch_message(455 downto 452);
 ch_message_align(1839 downto 1824) <= ch_message(459 downto 456) & ch_message(459 downto 456) & ch_message(459 downto 456) & ch_message(459 downto 456);
 ch_message_align(1855 downto 1840) <= ch_message(463 downto 460) & ch_message(463 downto 460) & ch_message(463 downto 460) & ch_message(463 downto 460);
 ch_message_align(1871 downto 1856) <= ch_message(467 downto 464) & ch_message(467 downto 464) & ch_message(467 downto 464) & ch_message(467 downto 464);
 ch_message_align(1887 downto 1872) <= ch_message(471 downto 468) & ch_message(471 downto 468) & ch_message(471 downto 468) & ch_message(471 downto 468);
 ch_message_align(1903 downto 1888) <= ch_message(475 downto 472) & ch_message(475 downto 472) & ch_message(475 downto 472) & ch_message(475 downto 472);
 ch_message_align(1919 downto 1904) <= ch_message(479 downto 476) & ch_message(479 downto 476) & ch_message(479 downto 476) & ch_message(479 downto 476);
 ch_message_align(1935 downto 1920) <= ch_message(483 downto 480) & ch_message(483 downto 480) & ch_message(483 downto 480) & ch_message(483 downto 480);
 ch_message_align(1951 downto 1936) <= ch_message(487 downto 484) & ch_message(487 downto 484) & ch_message(487 downto 484) & ch_message(487 downto 484);
 ch_message_align(1967 downto 1952) <= ch_message(491 downto 488) & ch_message(491 downto 488) & ch_message(491 downto 488) & ch_message(491 downto 488);
 ch_message_align(1983 downto 1968) <= ch_message(495 downto 492) & ch_message(495 downto 492) & ch_message(495 downto 492) & ch_message(495 downto 492);
 ch_message_align(1999 downto 1984) <= ch_message(499 downto 496) & ch_message(499 downto 496) & ch_message(499 downto 496) & ch_message(499 downto 496);
 ch_message_align(2015 downto 2000) <= ch_message(503 downto 500) & ch_message(503 downto 500) & ch_message(503 downto 500) & ch_message(503 downto 500);
 ch_message_align(2031 downto 2016) <= ch_message(507 downto 504) & ch_message(507 downto 504) & ch_message(507 downto 504) & ch_message(507 downto 504);
 ch_message_align(2047 downto 2032) <= ch_message(511 downto 508) & ch_message(511 downto 508) & ch_message(511 downto 508) & ch_message(511 downto 508);


   v_message_align(3 downto 0)<=ch_message_align(3 downto 0) when (mux_control='1') else v_message(3 downto 0);
   v_message_align(7 downto 4)<=ch_message_align(19 downto 16) when (mux_control='1') else v_message(19 downto 16);
   v_message_align(11 downto 8)<=ch_message_align(35 downto 32) when (mux_control='1') else v_message(35 downto 32);
   v_message_align(15 downto 12)<=ch_message_align(51 downto 48) when (mux_control='1') else v_message(51 downto 48);
   v_message_align(19 downto 16)<=ch_message_align(67 downto 64) when (mux_control='1') else v_message(67 downto 64);
   v_message_align(23 downto 20)<=ch_message_align(83 downto 80) when (mux_control='1') else v_message(83 downto 80);
   v_message_align(27 downto 24)<=ch_message_align(99 downto 96) when (mux_control='1') else v_message(99 downto 96);
   v_message_align(31 downto 28)<=ch_message_align(115 downto 112) when (mux_control='1') else v_message(115 downto 112);
   v_message_align(35 downto 32)<=ch_message_align(131 downto 128) when (mux_control='1') else v_message(131 downto 128);
   v_message_align(39 downto 36)<=ch_message_align(147 downto 144) when (mux_control='1') else v_message(147 downto 144);
   v_message_align(43 downto 40)<=ch_message_align(163 downto 160) when (mux_control='1') else v_message(163 downto 160);
   v_message_align(47 downto 44)<=ch_message_align(179 downto 176) when (mux_control='1') else v_message(179 downto 176);
   v_message_align(51 downto 48)<=ch_message_align(195 downto 192) when (mux_control='1') else v_message(195 downto 192);
   v_message_align(55 downto 52)<=ch_message_align(211 downto 208) when (mux_control='1') else v_message(211 downto 208);
   v_message_align(59 downto 56)<=ch_message_align(227 downto 224) when (mux_control='1') else v_message(227 downto 224);
   v_message_align(63 downto 60)<=ch_message_align(243 downto 240) when (mux_control='1') else v_message(243 downto 240);
   v_message_align(67 downto 64)<=ch_message_align(259 downto 256) when (mux_control='1') else v_message(259 downto 256);
   v_message_align(71 downto 68)<=ch_message_align(275 downto 272) when (mux_control='1') else v_message(275 downto 272);
   v_message_align(75 downto 72)<=ch_message_align(291 downto 288) when (mux_control='1') else v_message(291 downto 288);
   v_message_align(79 downto 76)<=ch_message_align(307 downto 304) when (mux_control='1') else v_message(307 downto 304);
   v_message_align(83 downto 80)<=ch_message_align(323 downto 320) when (mux_control='1') else v_message(323 downto 320);
   v_message_align(87 downto 84)<=ch_message_align(339 downto 336) when (mux_control='1') else v_message(339 downto 336);
   v_message_align(91 downto 88)<=ch_message_align(355 downto 352) when (mux_control='1') else v_message(355 downto 352);
   v_message_align(95 downto 92)<=ch_message_align(371 downto 368) when (mux_control='1') else v_message(371 downto 368);
   v_message_align(99 downto 96)<=ch_message_align(387 downto 384) when (mux_control='1') else v_message(387 downto 384);
   v_message_align(103 downto 100)<=ch_message_align(403 downto 400) when (mux_control='1') else v_message(403 downto 400);
   v_message_align(107 downto 104)<=ch_message_align(419 downto 416) when (mux_control='1') else v_message(419 downto 416);
   v_message_align(111 downto 108)<=ch_message_align(435 downto 432) when (mux_control='1') else v_message(435 downto 432);
   v_message_align(115 downto 112)<=ch_message_align(451 downto 448) when (mux_control='1') else v_message(451 downto 448);
   v_message_align(119 downto 116)<=ch_message_align(467 downto 464) when (mux_control='1') else v_message(467 downto 464);
   v_message_align(123 downto 120)<=ch_message_align(483 downto 480) when (mux_control='1') else v_message(483 downto 480);
   v_message_align(127 downto 124)<=ch_message_align(499 downto 496) when (mux_control='1') else v_message(499 downto 496);
   v_message_align(131 downto 128)<=ch_message_align(515 downto 512) when (mux_control='1') else v_message(515 downto 512);
   v_message_align(135 downto 132)<=ch_message_align(531 downto 528) when (mux_control='1') else v_message(531 downto 528);
   v_message_align(139 downto 136)<=ch_message_align(547 downto 544) when (mux_control='1') else v_message(547 downto 544);
   v_message_align(143 downto 140)<=ch_message_align(563 downto 560) when (mux_control='1') else v_message(563 downto 560);
   v_message_align(147 downto 144)<=ch_message_align(579 downto 576) when (mux_control='1') else v_message(579 downto 576);
   v_message_align(151 downto 148)<=ch_message_align(595 downto 592) when (mux_control='1') else v_message(595 downto 592);
   v_message_align(155 downto 152)<=ch_message_align(611 downto 608) when (mux_control='1') else v_message(611 downto 608);
   v_message_align(159 downto 156)<=ch_message_align(627 downto 624) when (mux_control='1') else v_message(627 downto 624);
   v_message_align(163 downto 160)<=ch_message_align(643 downto 640) when (mux_control='1') else v_message(643 downto 640);
   v_message_align(167 downto 164)<=ch_message_align(659 downto 656) when (mux_control='1') else v_message(659 downto 656);
   v_message_align(171 downto 168)<=ch_message_align(675 downto 672) when (mux_control='1') else v_message(675 downto 672);
   v_message_align(175 downto 172)<=ch_message_align(691 downto 688) when (mux_control='1') else v_message(691 downto 688);
   v_message_align(179 downto 176)<=ch_message_align(707 downto 704) when (mux_control='1') else v_message(707 downto 704);
   v_message_align(183 downto 180)<=ch_message_align(723 downto 720) when (mux_control='1') else v_message(723 downto 720);
   v_message_align(187 downto 184)<=ch_message_align(739 downto 736) when (mux_control='1') else v_message(739 downto 736);
   v_message_align(191 downto 188)<=ch_message_align(755 downto 752) when (mux_control='1') else v_message(755 downto 752);
   v_message_align(195 downto 192)<=ch_message_align(771 downto 768) when (mux_control='1') else v_message(771 downto 768);
   v_message_align(199 downto 196)<=ch_message_align(787 downto 784) when (mux_control='1') else v_message(787 downto 784);
   v_message_align(203 downto 200)<=ch_message_align(803 downto 800) when (mux_control='1') else v_message(803 downto 800);
   v_message_align(207 downto 204)<=ch_message_align(819 downto 816) when (mux_control='1') else v_message(819 downto 816);
   v_message_align(211 downto 208)<=ch_message_align(835 downto 832) when (mux_control='1') else v_message(835 downto 832);
   v_message_align(215 downto 212)<=ch_message_align(851 downto 848) when (mux_control='1') else v_message(851 downto 848);
   v_message_align(219 downto 216)<=ch_message_align(867 downto 864) when (mux_control='1') else v_message(867 downto 864);
   v_message_align(223 downto 220)<=ch_message_align(883 downto 880) when (mux_control='1') else v_message(883 downto 880);
   v_message_align(227 downto 224)<=ch_message_align(899 downto 896) when (mux_control='1') else v_message(899 downto 896);
   v_message_align(231 downto 228)<=ch_message_align(915 downto 912) when (mux_control='1') else v_message(915 downto 912);
   v_message_align(235 downto 232)<=ch_message_align(931 downto 928) when (mux_control='1') else v_message(931 downto 928);
   v_message_align(239 downto 236)<=ch_message_align(947 downto 944) when (mux_control='1') else v_message(947 downto 944);
   v_message_align(243 downto 240)<=ch_message_align(963 downto 960) when (mux_control='1') else v_message(963 downto 960);
   v_message_align(247 downto 244)<=ch_message_align(979 downto 976) when (mux_control='1') else v_message(979 downto 976);
   v_message_align(251 downto 248)<=ch_message_align(995 downto 992) when (mux_control='1') else v_message(995 downto 992);
   v_message_align(255 downto 252)<=ch_message_align(1011 downto 1008) when (mux_control='1') else v_message(1011 downto 1008);
   v_message_align(259 downto 256)<=ch_message_align(1027 downto 1024) when (mux_control='1') else v_message(1027 downto 1024);
   v_message_align(263 downto 260)<=ch_message_align(1043 downto 1040) when (mux_control='1') else v_message(1043 downto 1040);
   v_message_align(267 downto 264)<=ch_message_align(1059 downto 1056) when (mux_control='1') else v_message(1059 downto 1056);
   v_message_align(271 downto 268)<=ch_message_align(1075 downto 1072) when (mux_control='1') else v_message(1075 downto 1072);
   v_message_align(275 downto 272)<=ch_message_align(1091 downto 1088) when (mux_control='1') else v_message(1091 downto 1088);
   v_message_align(279 downto 276)<=ch_message_align(1107 downto 1104) when (mux_control='1') else v_message(1107 downto 1104);
   v_message_align(283 downto 280)<=ch_message_align(1123 downto 1120) when (mux_control='1') else v_message(1123 downto 1120);
   v_message_align(287 downto 284)<=ch_message_align(1139 downto 1136) when (mux_control='1') else v_message(1139 downto 1136);
   v_message_align(291 downto 288)<=ch_message_align(1155 downto 1152) when (mux_control='1') else v_message(1155 downto 1152);
   v_message_align(295 downto 292)<=ch_message_align(1171 downto 1168) when (mux_control='1') else v_message(1171 downto 1168);
   v_message_align(299 downto 296)<=ch_message_align(1187 downto 1184) when (mux_control='1') else v_message(1187 downto 1184);
   v_message_align(303 downto 300)<=ch_message_align(1203 downto 1200) when (mux_control='1') else v_message(1203 downto 1200);
   v_message_align(307 downto 304)<=ch_message_align(1219 downto 1216) when (mux_control='1') else v_message(1219 downto 1216);
   v_message_align(311 downto 308)<=ch_message_align(1235 downto 1232) when (mux_control='1') else v_message(1235 downto 1232);
   v_message_align(315 downto 312)<=ch_message_align(1251 downto 1248) when (mux_control='1') else v_message(1251 downto 1248);
   v_message_align(319 downto 316)<=ch_message_align(1267 downto 1264) when (mux_control='1') else v_message(1267 downto 1264);
   v_message_align(323 downto 320)<=ch_message_align(1283 downto 1280) when (mux_control='1') else v_message(1283 downto 1280);
   v_message_align(327 downto 324)<=ch_message_align(1299 downto 1296) when (mux_control='1') else v_message(1299 downto 1296);
   v_message_align(331 downto 328)<=ch_message_align(1315 downto 1312) when (mux_control='1') else v_message(1315 downto 1312);
   v_message_align(335 downto 332)<=ch_message_align(1331 downto 1328) when (mux_control='1') else v_message(1331 downto 1328);
   v_message_align(339 downto 336)<=ch_message_align(1347 downto 1344) when (mux_control='1') else v_message(1347 downto 1344);
   v_message_align(343 downto 340)<=ch_message_align(1363 downto 1360) when (mux_control='1') else v_message(1363 downto 1360);
   v_message_align(347 downto 344)<=ch_message_align(1379 downto 1376) when (mux_control='1') else v_message(1379 downto 1376);
   v_message_align(351 downto 348)<=ch_message_align(1395 downto 1392) when (mux_control='1') else v_message(1395 downto 1392);
   v_message_align(355 downto 352)<=ch_message_align(1411 downto 1408) when (mux_control='1') else v_message(1411 downto 1408);
   v_message_align(359 downto 356)<=ch_message_align(1427 downto 1424) when (mux_control='1') else v_message(1427 downto 1424);
   v_message_align(363 downto 360)<=ch_message_align(1443 downto 1440) when (mux_control='1') else v_message(1443 downto 1440);
   v_message_align(367 downto 364)<=ch_message_align(1459 downto 1456) when (mux_control='1') else v_message(1459 downto 1456);
   v_message_align(371 downto 368)<=ch_message_align(1475 downto 1472) when (mux_control='1') else v_message(1475 downto 1472);
   v_message_align(375 downto 372)<=ch_message_align(1491 downto 1488) when (mux_control='1') else v_message(1491 downto 1488);
   v_message_align(379 downto 376)<=ch_message_align(1507 downto 1504) when (mux_control='1') else v_message(1507 downto 1504);
   v_message_align(383 downto 380)<=ch_message_align(1523 downto 1520) when (mux_control='1') else v_message(1523 downto 1520);
   v_message_align(387 downto 384)<=ch_message_align(1539 downto 1536) when (mux_control='1') else v_message(1539 downto 1536);
   v_message_align(391 downto 388)<=ch_message_align(1555 downto 1552) when (mux_control='1') else v_message(1555 downto 1552);
   v_message_align(395 downto 392)<=ch_message_align(1571 downto 1568) when (mux_control='1') else v_message(1571 downto 1568);
   v_message_align(399 downto 396)<=ch_message_align(1587 downto 1584) when (mux_control='1') else v_message(1587 downto 1584);
   v_message_align(403 downto 400)<=ch_message_align(1603 downto 1600) when (mux_control='1') else v_message(1603 downto 1600);
   v_message_align(407 downto 404)<=ch_message_align(1619 downto 1616) when (mux_control='1') else v_message(1619 downto 1616);
   v_message_align(411 downto 408)<=ch_message_align(1635 downto 1632) when (mux_control='1') else v_message(1635 downto 1632);
   v_message_align(415 downto 412)<=ch_message_align(1651 downto 1648) when (mux_control='1') else v_message(1651 downto 1648);
   v_message_align(419 downto 416)<=ch_message_align(1667 downto 1664) when (mux_control='1') else v_message(1667 downto 1664);
   v_message_align(423 downto 420)<=ch_message_align(1683 downto 1680) when (mux_control='1') else v_message(1683 downto 1680);
   v_message_align(427 downto 424)<=ch_message_align(1699 downto 1696) when (mux_control='1') else v_message(1699 downto 1696);
   v_message_align(431 downto 428)<=ch_message_align(1715 downto 1712) when (mux_control='1') else v_message(1715 downto 1712);
   v_message_align(435 downto 432)<=ch_message_align(1731 downto 1728) when (mux_control='1') else v_message(1731 downto 1728);
   v_message_align(439 downto 436)<=ch_message_align(1747 downto 1744) when (mux_control='1') else v_message(1747 downto 1744);
   v_message_align(443 downto 440)<=ch_message_align(1763 downto 1760) when (mux_control='1') else v_message(1763 downto 1760);
   v_message_align(447 downto 444)<=ch_message_align(1779 downto 1776) when (mux_control='1') else v_message(1779 downto 1776);
   v_message_align(451 downto 448)<=ch_message_align(1795 downto 1792) when (mux_control='1') else v_message(1795 downto 1792);
   v_message_align(455 downto 452)<=ch_message_align(1811 downto 1808) when (mux_control='1') else v_message(1811 downto 1808);
   v_message_align(459 downto 456)<=ch_message_align(1827 downto 1824) when (mux_control='1') else v_message(1827 downto 1824);
   v_message_align(463 downto 460)<=ch_message_align(1843 downto 1840) when (mux_control='1') else v_message(1843 downto 1840);
   v_message_align(467 downto 464)<=ch_message_align(1859 downto 1856) when (mux_control='1') else v_message(1859 downto 1856);
   v_message_align(471 downto 468)<=ch_message_align(1875 downto 1872) when (mux_control='1') else v_message(1875 downto 1872);
   v_message_align(475 downto 472)<=ch_message_align(1891 downto 1888) when (mux_control='1') else v_message(1891 downto 1888);
   v_message_align(479 downto 476)<=ch_message_align(1907 downto 1904) when (mux_control='1') else v_message(1907 downto 1904);
   v_message_align(483 downto 480)<=ch_message_align(1923 downto 1920) when (mux_control='1') else v_message(1923 downto 1920);
   v_message_align(487 downto 484)<=ch_message_align(1939 downto 1936) when (mux_control='1') else v_message(1939 downto 1936);
   v_message_align(491 downto 488)<=ch_message_align(1955 downto 1952) when (mux_control='1') else v_message(1955 downto 1952);
   v_message_align(495 downto 492)<=ch_message_align(1971 downto 1968) when (mux_control='1') else v_message(1971 downto 1968);
   v_message_align(499 downto 496)<=ch_message_align(1987 downto 1984) when (mux_control='1') else v_message(1987 downto 1984);
   v_message_align(503 downto 500)<=ch_message_align(2003 downto 2000) when (mux_control='1') else v_message(2003 downto 2000);
   v_message_align(507 downto 504)<=ch_message_align(2019 downto 2016) when (mux_control='1') else v_message(2019 downto 2016);
   v_message_align(511 downto 508)<=ch_message_align(2035 downto 2032) when (mux_control='1') else v_message(2035 downto 2032);
   v_message_align(515 downto 512)<=ch_message_align(11 downto 8) when (mux_control='1') else v_message(11 downto 8);
   v_message_align(519 downto 516)<=ch_message_align(27 downto 24) when (mux_control='1') else v_message(27 downto 24);
   v_message_align(523 downto 520)<=ch_message_align(43 downto 40) when (mux_control='1') else v_message(43 downto 40);
   v_message_align(527 downto 524)<=ch_message_align(59 downto 56) when (mux_control='1') else v_message(59 downto 56);
   v_message_align(531 downto 528)<=ch_message_align(75 downto 72) when (mux_control='1') else v_message(75 downto 72);
   v_message_align(535 downto 532)<=ch_message_align(91 downto 88) when (mux_control='1') else v_message(91 downto 88);
   v_message_align(539 downto 536)<=ch_message_align(107 downto 104) when (mux_control='1') else v_message(107 downto 104);
   v_message_align(543 downto 540)<=ch_message_align(123 downto 120) when (mux_control='1') else v_message(123 downto 120);
   v_message_align(547 downto 544)<=ch_message_align(139 downto 136) when (mux_control='1') else v_message(139 downto 136);
   v_message_align(551 downto 548)<=ch_message_align(155 downto 152) when (mux_control='1') else v_message(155 downto 152);
   v_message_align(555 downto 552)<=ch_message_align(171 downto 168) when (mux_control='1') else v_message(171 downto 168);
   v_message_align(559 downto 556)<=ch_message_align(187 downto 184) when (mux_control='1') else v_message(187 downto 184);
   v_message_align(563 downto 560)<=ch_message_align(203 downto 200) when (mux_control='1') else v_message(203 downto 200);
   v_message_align(567 downto 564)<=ch_message_align(219 downto 216) when (mux_control='1') else v_message(219 downto 216);
   v_message_align(571 downto 568)<=ch_message_align(235 downto 232) when (mux_control='1') else v_message(235 downto 232);
   v_message_align(575 downto 572)<=ch_message_align(251 downto 248) when (mux_control='1') else v_message(251 downto 248);
   v_message_align(579 downto 576)<=ch_message_align(267 downto 264) when (mux_control='1') else v_message(267 downto 264);
   v_message_align(583 downto 580)<=ch_message_align(283 downto 280) when (mux_control='1') else v_message(283 downto 280);
   v_message_align(587 downto 584)<=ch_message_align(299 downto 296) when (mux_control='1') else v_message(299 downto 296);
   v_message_align(591 downto 588)<=ch_message_align(315 downto 312) when (mux_control='1') else v_message(315 downto 312);
   v_message_align(595 downto 592)<=ch_message_align(331 downto 328) when (mux_control='1') else v_message(331 downto 328);
   v_message_align(599 downto 596)<=ch_message_align(347 downto 344) when (mux_control='1') else v_message(347 downto 344);
   v_message_align(603 downto 600)<=ch_message_align(363 downto 360) when (mux_control='1') else v_message(363 downto 360);
   v_message_align(607 downto 604)<=ch_message_align(379 downto 376) when (mux_control='1') else v_message(379 downto 376);
   v_message_align(611 downto 608)<=ch_message_align(395 downto 392) when (mux_control='1') else v_message(395 downto 392);
   v_message_align(615 downto 612)<=ch_message_align(411 downto 408) when (mux_control='1') else v_message(411 downto 408);
   v_message_align(619 downto 616)<=ch_message_align(427 downto 424) when (mux_control='1') else v_message(427 downto 424);
   v_message_align(623 downto 620)<=ch_message_align(443 downto 440) when (mux_control='1') else v_message(443 downto 440);
   v_message_align(627 downto 624)<=ch_message_align(459 downto 456) when (mux_control='1') else v_message(459 downto 456);
   v_message_align(631 downto 628)<=ch_message_align(475 downto 472) when (mux_control='1') else v_message(475 downto 472);
   v_message_align(635 downto 632)<=ch_message_align(491 downto 488) when (mux_control='1') else v_message(491 downto 488);
   v_message_align(639 downto 636)<=ch_message_align(507 downto 504) when (mux_control='1') else v_message(507 downto 504);
   v_message_align(643 downto 640)<=ch_message_align(523 downto 520) when (mux_control='1') else v_message(523 downto 520);
   v_message_align(647 downto 644)<=ch_message_align(539 downto 536) when (mux_control='1') else v_message(539 downto 536);
   v_message_align(651 downto 648)<=ch_message_align(555 downto 552) when (mux_control='1') else v_message(555 downto 552);
   v_message_align(655 downto 652)<=ch_message_align(571 downto 568) when (mux_control='1') else v_message(571 downto 568);
   v_message_align(659 downto 656)<=ch_message_align(587 downto 584) when (mux_control='1') else v_message(587 downto 584);
   v_message_align(663 downto 660)<=ch_message_align(603 downto 600) when (mux_control='1') else v_message(603 downto 600);
   v_message_align(667 downto 664)<=ch_message_align(619 downto 616) when (mux_control='1') else v_message(619 downto 616);
   v_message_align(671 downto 668)<=ch_message_align(635 downto 632) when (mux_control='1') else v_message(635 downto 632);
   v_message_align(675 downto 672)<=ch_message_align(651 downto 648) when (mux_control='1') else v_message(651 downto 648);
   v_message_align(679 downto 676)<=ch_message_align(667 downto 664) when (mux_control='1') else v_message(667 downto 664);
   v_message_align(683 downto 680)<=ch_message_align(683 downto 680) when (mux_control='1') else v_message(683 downto 680);
   v_message_align(687 downto 684)<=ch_message_align(699 downto 696) when (mux_control='1') else v_message(699 downto 696);
   v_message_align(691 downto 688)<=ch_message_align(715 downto 712) when (mux_control='1') else v_message(715 downto 712);
   v_message_align(695 downto 692)<=ch_message_align(731 downto 728) when (mux_control='1') else v_message(731 downto 728);
   v_message_align(699 downto 696)<=ch_message_align(747 downto 744) when (mux_control='1') else v_message(747 downto 744);
   v_message_align(703 downto 700)<=ch_message_align(763 downto 760) when (mux_control='1') else v_message(763 downto 760);
   v_message_align(707 downto 704)<=ch_message_align(779 downto 776) when (mux_control='1') else v_message(779 downto 776);
   v_message_align(711 downto 708)<=ch_message_align(795 downto 792) when (mux_control='1') else v_message(795 downto 792);
   v_message_align(715 downto 712)<=ch_message_align(811 downto 808) when (mux_control='1') else v_message(811 downto 808);
   v_message_align(719 downto 716)<=ch_message_align(827 downto 824) when (mux_control='1') else v_message(827 downto 824);
   v_message_align(723 downto 720)<=ch_message_align(843 downto 840) when (mux_control='1') else v_message(843 downto 840);
   v_message_align(727 downto 724)<=ch_message_align(859 downto 856) when (mux_control='1') else v_message(859 downto 856);
   v_message_align(731 downto 728)<=ch_message_align(875 downto 872) when (mux_control='1') else v_message(875 downto 872);
   v_message_align(735 downto 732)<=ch_message_align(891 downto 888) when (mux_control='1') else v_message(891 downto 888);
   v_message_align(739 downto 736)<=ch_message_align(907 downto 904) when (mux_control='1') else v_message(907 downto 904);
   v_message_align(743 downto 740)<=ch_message_align(923 downto 920) when (mux_control='1') else v_message(923 downto 920);
   v_message_align(747 downto 744)<=ch_message_align(939 downto 936) when (mux_control='1') else v_message(939 downto 936);
   v_message_align(751 downto 748)<=ch_message_align(955 downto 952) when (mux_control='1') else v_message(955 downto 952);
   v_message_align(755 downto 752)<=ch_message_align(971 downto 968) when (mux_control='1') else v_message(971 downto 968);
   v_message_align(759 downto 756)<=ch_message_align(987 downto 984) when (mux_control='1') else v_message(987 downto 984);
   v_message_align(763 downto 760)<=ch_message_align(1003 downto 1000) when (mux_control='1') else v_message(1003 downto 1000);
   v_message_align(767 downto 764)<=ch_message_align(1019 downto 1016) when (mux_control='1') else v_message(1019 downto 1016);
   v_message_align(771 downto 768)<=ch_message_align(1035 downto 1032) when (mux_control='1') else v_message(1035 downto 1032);
   v_message_align(775 downto 772)<=ch_message_align(1051 downto 1048) when (mux_control='1') else v_message(1051 downto 1048);
   v_message_align(779 downto 776)<=ch_message_align(1067 downto 1064) when (mux_control='1') else v_message(1067 downto 1064);
   v_message_align(783 downto 780)<=ch_message_align(1083 downto 1080) when (mux_control='1') else v_message(1083 downto 1080);
   v_message_align(787 downto 784)<=ch_message_align(1099 downto 1096) when (mux_control='1') else v_message(1099 downto 1096);
   v_message_align(791 downto 788)<=ch_message_align(1115 downto 1112) when (mux_control='1') else v_message(1115 downto 1112);
   v_message_align(795 downto 792)<=ch_message_align(1131 downto 1128) when (mux_control='1') else v_message(1131 downto 1128);
   v_message_align(799 downto 796)<=ch_message_align(1147 downto 1144) when (mux_control='1') else v_message(1147 downto 1144);
   v_message_align(803 downto 800)<=ch_message_align(1163 downto 1160) when (mux_control='1') else v_message(1163 downto 1160);
   v_message_align(807 downto 804)<=ch_message_align(1179 downto 1176) when (mux_control='1') else v_message(1179 downto 1176);
   v_message_align(811 downto 808)<=ch_message_align(1195 downto 1192) when (mux_control='1') else v_message(1195 downto 1192);
   v_message_align(815 downto 812)<=ch_message_align(1211 downto 1208) when (mux_control='1') else v_message(1211 downto 1208);
   v_message_align(819 downto 816)<=ch_message_align(1227 downto 1224) when (mux_control='1') else v_message(1227 downto 1224);
   v_message_align(823 downto 820)<=ch_message_align(1243 downto 1240) when (mux_control='1') else v_message(1243 downto 1240);
   v_message_align(827 downto 824)<=ch_message_align(1259 downto 1256) when (mux_control='1') else v_message(1259 downto 1256);
   v_message_align(831 downto 828)<=ch_message_align(1275 downto 1272) when (mux_control='1') else v_message(1275 downto 1272);
   v_message_align(835 downto 832)<=ch_message_align(1291 downto 1288) when (mux_control='1') else v_message(1291 downto 1288);
   v_message_align(839 downto 836)<=ch_message_align(1307 downto 1304) when (mux_control='1') else v_message(1307 downto 1304);
   v_message_align(843 downto 840)<=ch_message_align(1323 downto 1320) when (mux_control='1') else v_message(1323 downto 1320);
   v_message_align(847 downto 844)<=ch_message_align(1339 downto 1336) when (mux_control='1') else v_message(1339 downto 1336);
   v_message_align(851 downto 848)<=ch_message_align(1355 downto 1352) when (mux_control='1') else v_message(1355 downto 1352);
   v_message_align(855 downto 852)<=ch_message_align(1371 downto 1368) when (mux_control='1') else v_message(1371 downto 1368);
   v_message_align(859 downto 856)<=ch_message_align(1387 downto 1384) when (mux_control='1') else v_message(1387 downto 1384);
   v_message_align(863 downto 860)<=ch_message_align(1403 downto 1400) when (mux_control='1') else v_message(1403 downto 1400);
   v_message_align(867 downto 864)<=ch_message_align(1419 downto 1416) when (mux_control='1') else v_message(1419 downto 1416);
   v_message_align(871 downto 868)<=ch_message_align(1435 downto 1432) when (mux_control='1') else v_message(1435 downto 1432);
   v_message_align(875 downto 872)<=ch_message_align(1451 downto 1448) when (mux_control='1') else v_message(1451 downto 1448);
   v_message_align(879 downto 876)<=ch_message_align(1467 downto 1464) when (mux_control='1') else v_message(1467 downto 1464);
   v_message_align(883 downto 880)<=ch_message_align(1483 downto 1480) when (mux_control='1') else v_message(1483 downto 1480);
   v_message_align(887 downto 884)<=ch_message_align(1499 downto 1496) when (mux_control='1') else v_message(1499 downto 1496);
   v_message_align(891 downto 888)<=ch_message_align(1515 downto 1512) when (mux_control='1') else v_message(1515 downto 1512);
   v_message_align(895 downto 892)<=ch_message_align(1531 downto 1528) when (mux_control='1') else v_message(1531 downto 1528);
   v_message_align(899 downto 896)<=ch_message_align(1547 downto 1544) when (mux_control='1') else v_message(1547 downto 1544);
   v_message_align(903 downto 900)<=ch_message_align(1563 downto 1560) when (mux_control='1') else v_message(1563 downto 1560);
   v_message_align(907 downto 904)<=ch_message_align(1579 downto 1576) when (mux_control='1') else v_message(1579 downto 1576);
   v_message_align(911 downto 908)<=ch_message_align(1595 downto 1592) when (mux_control='1') else v_message(1595 downto 1592);
   v_message_align(915 downto 912)<=ch_message_align(1611 downto 1608) when (mux_control='1') else v_message(1611 downto 1608);
   v_message_align(919 downto 916)<=ch_message_align(1627 downto 1624) when (mux_control='1') else v_message(1627 downto 1624);
   v_message_align(923 downto 920)<=ch_message_align(1643 downto 1640) when (mux_control='1') else v_message(1643 downto 1640);
   v_message_align(927 downto 924)<=ch_message_align(1659 downto 1656) when (mux_control='1') else v_message(1659 downto 1656);
   v_message_align(931 downto 928)<=ch_message_align(1675 downto 1672) when (mux_control='1') else v_message(1675 downto 1672);
   v_message_align(935 downto 932)<=ch_message_align(1691 downto 1688) when (mux_control='1') else v_message(1691 downto 1688);
   v_message_align(939 downto 936)<=ch_message_align(1707 downto 1704) when (mux_control='1') else v_message(1707 downto 1704);
   v_message_align(943 downto 940)<=ch_message_align(1723 downto 1720) when (mux_control='1') else v_message(1723 downto 1720);
   v_message_align(947 downto 944)<=ch_message_align(1739 downto 1736) when (mux_control='1') else v_message(1739 downto 1736);
   v_message_align(951 downto 948)<=ch_message_align(1755 downto 1752) when (mux_control='1') else v_message(1755 downto 1752);
   v_message_align(955 downto 952)<=ch_message_align(1771 downto 1768) when (mux_control='1') else v_message(1771 downto 1768);
   v_message_align(959 downto 956)<=ch_message_align(1787 downto 1784) when (mux_control='1') else v_message(1787 downto 1784);
   v_message_align(963 downto 960)<=ch_message_align(1803 downto 1800) when (mux_control='1') else v_message(1803 downto 1800);
   v_message_align(967 downto 964)<=ch_message_align(1819 downto 1816) when (mux_control='1') else v_message(1819 downto 1816);
   v_message_align(971 downto 968)<=ch_message_align(1835 downto 1832) when (mux_control='1') else v_message(1835 downto 1832);
   v_message_align(975 downto 972)<=ch_message_align(1851 downto 1848) when (mux_control='1') else v_message(1851 downto 1848);
   v_message_align(979 downto 976)<=ch_message_align(1867 downto 1864) when (mux_control='1') else v_message(1867 downto 1864);
   v_message_align(983 downto 980)<=ch_message_align(1883 downto 1880) when (mux_control='1') else v_message(1883 downto 1880);
   v_message_align(987 downto 984)<=ch_message_align(1899 downto 1896) when (mux_control='1') else v_message(1899 downto 1896);
   v_message_align(991 downto 988)<=ch_message_align(1915 downto 1912) when (mux_control='1') else v_message(1915 downto 1912);
   v_message_align(995 downto 992)<=ch_message_align(1931 downto 1928) when (mux_control='1') else v_message(1931 downto 1928);
   v_message_align(999 downto 996)<=ch_message_align(1947 downto 1944) when (mux_control='1') else v_message(1947 downto 1944);
   v_message_align(1003 downto 1000)<=ch_message_align(1963 downto 1960) when (mux_control='1') else v_message(1963 downto 1960);
   v_message_align(1007 downto 1004)<=ch_message_align(1979 downto 1976) when (mux_control='1') else v_message(1979 downto 1976);
   v_message_align(1011 downto 1008)<=ch_message_align(1995 downto 1992) when (mux_control='1') else v_message(1995 downto 1992);
   v_message_align(1015 downto 1012)<=ch_message_align(2011 downto 2008) when (mux_control='1') else v_message(2011 downto 2008);
   v_message_align(1019 downto 1016)<=ch_message_align(2027 downto 2024) when (mux_control='1') else v_message(2027 downto 2024);
   v_message_align(1023 downto 1020)<=ch_message_align(2043 downto 2040) when (mux_control='1') else v_message(2043 downto 2040);
   v_message_align(1027 downto 1024)<=ch_message_align(7 downto 4) when (mux_control='1') else v_message(7 downto 4);
   v_message_align(1031 downto 1028)<=ch_message_align(23 downto 20) when (mux_control='1') else v_message(23 downto 20);
   v_message_align(1035 downto 1032)<=ch_message_align(39 downto 36) when (mux_control='1') else v_message(39 downto 36);
   v_message_align(1039 downto 1036)<=ch_message_align(55 downto 52) when (mux_control='1') else v_message(55 downto 52);
   v_message_align(1043 downto 1040)<=ch_message_align(71 downto 68) when (mux_control='1') else v_message(71 downto 68);
   v_message_align(1047 downto 1044)<=ch_message_align(87 downto 84) when (mux_control='1') else v_message(87 downto 84);
   v_message_align(1051 downto 1048)<=ch_message_align(103 downto 100) when (mux_control='1') else v_message(103 downto 100);
   v_message_align(1055 downto 1052)<=ch_message_align(119 downto 116) when (mux_control='1') else v_message(119 downto 116);
   v_message_align(1059 downto 1056)<=ch_message_align(135 downto 132) when (mux_control='1') else v_message(135 downto 132);
   v_message_align(1063 downto 1060)<=ch_message_align(151 downto 148) when (mux_control='1') else v_message(151 downto 148);
   v_message_align(1067 downto 1064)<=ch_message_align(167 downto 164) when (mux_control='1') else v_message(167 downto 164);
   v_message_align(1071 downto 1068)<=ch_message_align(183 downto 180) when (mux_control='1') else v_message(183 downto 180);
   v_message_align(1075 downto 1072)<=ch_message_align(199 downto 196) when (mux_control='1') else v_message(199 downto 196);
   v_message_align(1079 downto 1076)<=ch_message_align(215 downto 212) when (mux_control='1') else v_message(215 downto 212);
   v_message_align(1083 downto 1080)<=ch_message_align(231 downto 228) when (mux_control='1') else v_message(231 downto 228);
   v_message_align(1087 downto 1084)<=ch_message_align(247 downto 244) when (mux_control='1') else v_message(247 downto 244);
   v_message_align(1091 downto 1088)<=ch_message_align(263 downto 260) when (mux_control='1') else v_message(263 downto 260);
   v_message_align(1095 downto 1092)<=ch_message_align(279 downto 276) when (mux_control='1') else v_message(279 downto 276);
   v_message_align(1099 downto 1096)<=ch_message_align(295 downto 292) when (mux_control='1') else v_message(295 downto 292);
   v_message_align(1103 downto 1100)<=ch_message_align(311 downto 308) when (mux_control='1') else v_message(311 downto 308);
   v_message_align(1107 downto 1104)<=ch_message_align(327 downto 324) when (mux_control='1') else v_message(327 downto 324);
   v_message_align(1111 downto 1108)<=ch_message_align(343 downto 340) when (mux_control='1') else v_message(343 downto 340);
   v_message_align(1115 downto 1112)<=ch_message_align(359 downto 356) when (mux_control='1') else v_message(359 downto 356);
   v_message_align(1119 downto 1116)<=ch_message_align(375 downto 372) when (mux_control='1') else v_message(375 downto 372);
   v_message_align(1123 downto 1120)<=ch_message_align(391 downto 388) when (mux_control='1') else v_message(391 downto 388);
   v_message_align(1127 downto 1124)<=ch_message_align(407 downto 404) when (mux_control='1') else v_message(407 downto 404);
   v_message_align(1131 downto 1128)<=ch_message_align(423 downto 420) when (mux_control='1') else v_message(423 downto 420);
   v_message_align(1135 downto 1132)<=ch_message_align(439 downto 436) when (mux_control='1') else v_message(439 downto 436);
   v_message_align(1139 downto 1136)<=ch_message_align(455 downto 452) when (mux_control='1') else v_message(455 downto 452);
   v_message_align(1143 downto 1140)<=ch_message_align(471 downto 468) when (mux_control='1') else v_message(471 downto 468);
   v_message_align(1147 downto 1144)<=ch_message_align(487 downto 484) when (mux_control='1') else v_message(487 downto 484);
   v_message_align(1151 downto 1148)<=ch_message_align(503 downto 500) when (mux_control='1') else v_message(503 downto 500);
   v_message_align(1155 downto 1152)<=ch_message_align(519 downto 516) when (mux_control='1') else v_message(519 downto 516);
   v_message_align(1159 downto 1156)<=ch_message_align(535 downto 532) when (mux_control='1') else v_message(535 downto 532);
   v_message_align(1163 downto 1160)<=ch_message_align(551 downto 548) when (mux_control='1') else v_message(551 downto 548);
   v_message_align(1167 downto 1164)<=ch_message_align(567 downto 564) when (mux_control='1') else v_message(567 downto 564);
   v_message_align(1171 downto 1168)<=ch_message_align(583 downto 580) when (mux_control='1') else v_message(583 downto 580);
   v_message_align(1175 downto 1172)<=ch_message_align(599 downto 596) when (mux_control='1') else v_message(599 downto 596);
   v_message_align(1179 downto 1176)<=ch_message_align(615 downto 612) when (mux_control='1') else v_message(615 downto 612);
   v_message_align(1183 downto 1180)<=ch_message_align(631 downto 628) when (mux_control='1') else v_message(631 downto 628);
   v_message_align(1187 downto 1184)<=ch_message_align(647 downto 644) when (mux_control='1') else v_message(647 downto 644);
   v_message_align(1191 downto 1188)<=ch_message_align(663 downto 660) when (mux_control='1') else v_message(663 downto 660);
   v_message_align(1195 downto 1192)<=ch_message_align(679 downto 676) when (mux_control='1') else v_message(679 downto 676);
   v_message_align(1199 downto 1196)<=ch_message_align(695 downto 692) when (mux_control='1') else v_message(695 downto 692);
   v_message_align(1203 downto 1200)<=ch_message_align(711 downto 708) when (mux_control='1') else v_message(711 downto 708);
   v_message_align(1207 downto 1204)<=ch_message_align(727 downto 724) when (mux_control='1') else v_message(727 downto 724);
   v_message_align(1211 downto 1208)<=ch_message_align(743 downto 740) when (mux_control='1') else v_message(743 downto 740);
   v_message_align(1215 downto 1212)<=ch_message_align(759 downto 756) when (mux_control='1') else v_message(759 downto 756);
   v_message_align(1219 downto 1216)<=ch_message_align(775 downto 772) when (mux_control='1') else v_message(775 downto 772);
   v_message_align(1223 downto 1220)<=ch_message_align(791 downto 788) when (mux_control='1') else v_message(791 downto 788);
   v_message_align(1227 downto 1224)<=ch_message_align(807 downto 804) when (mux_control='1') else v_message(807 downto 804);
   v_message_align(1231 downto 1228)<=ch_message_align(823 downto 820) when (mux_control='1') else v_message(823 downto 820);
   v_message_align(1235 downto 1232)<=ch_message_align(839 downto 836) when (mux_control='1') else v_message(839 downto 836);
   v_message_align(1239 downto 1236)<=ch_message_align(855 downto 852) when (mux_control='1') else v_message(855 downto 852);
   v_message_align(1243 downto 1240)<=ch_message_align(871 downto 868) when (mux_control='1') else v_message(871 downto 868);
   v_message_align(1247 downto 1244)<=ch_message_align(887 downto 884) when (mux_control='1') else v_message(887 downto 884);
   v_message_align(1251 downto 1248)<=ch_message_align(903 downto 900) when (mux_control='1') else v_message(903 downto 900);
   v_message_align(1255 downto 1252)<=ch_message_align(919 downto 916) when (mux_control='1') else v_message(919 downto 916);
   v_message_align(1259 downto 1256)<=ch_message_align(935 downto 932) when (mux_control='1') else v_message(935 downto 932);
   v_message_align(1263 downto 1260)<=ch_message_align(951 downto 948) when (mux_control='1') else v_message(951 downto 948);
   v_message_align(1267 downto 1264)<=ch_message_align(967 downto 964) when (mux_control='1') else v_message(967 downto 964);
   v_message_align(1271 downto 1268)<=ch_message_align(983 downto 980) when (mux_control='1') else v_message(983 downto 980);
   v_message_align(1275 downto 1272)<=ch_message_align(999 downto 996) when (mux_control='1') else v_message(999 downto 996);
   v_message_align(1279 downto 1276)<=ch_message_align(1015 downto 1012) when (mux_control='1') else v_message(1015 downto 1012);
   v_message_align(1283 downto 1280)<=ch_message_align(1031 downto 1028) when (mux_control='1') else v_message(1031 downto 1028);
   v_message_align(1287 downto 1284)<=ch_message_align(1047 downto 1044) when (mux_control='1') else v_message(1047 downto 1044);
   v_message_align(1291 downto 1288)<=ch_message_align(1063 downto 1060) when (mux_control='1') else v_message(1063 downto 1060);
   v_message_align(1295 downto 1292)<=ch_message_align(1079 downto 1076) when (mux_control='1') else v_message(1079 downto 1076);
   v_message_align(1299 downto 1296)<=ch_message_align(1095 downto 1092) when (mux_control='1') else v_message(1095 downto 1092);
   v_message_align(1303 downto 1300)<=ch_message_align(1111 downto 1108) when (mux_control='1') else v_message(1111 downto 1108);
   v_message_align(1307 downto 1304)<=ch_message_align(1127 downto 1124) when (mux_control='1') else v_message(1127 downto 1124);
   v_message_align(1311 downto 1308)<=ch_message_align(1143 downto 1140) when (mux_control='1') else v_message(1143 downto 1140);
   v_message_align(1315 downto 1312)<=ch_message_align(1159 downto 1156) when (mux_control='1') else v_message(1159 downto 1156);
   v_message_align(1319 downto 1316)<=ch_message_align(1175 downto 1172) when (mux_control='1') else v_message(1175 downto 1172);
   v_message_align(1323 downto 1320)<=ch_message_align(1191 downto 1188) when (mux_control='1') else v_message(1191 downto 1188);
   v_message_align(1327 downto 1324)<=ch_message_align(1207 downto 1204) when (mux_control='1') else v_message(1207 downto 1204);
   v_message_align(1331 downto 1328)<=ch_message_align(1223 downto 1220) when (mux_control='1') else v_message(1223 downto 1220);
   v_message_align(1335 downto 1332)<=ch_message_align(1239 downto 1236) when (mux_control='1') else v_message(1239 downto 1236);
   v_message_align(1339 downto 1336)<=ch_message_align(1255 downto 1252) when (mux_control='1') else v_message(1255 downto 1252);
   v_message_align(1343 downto 1340)<=ch_message_align(1271 downto 1268) when (mux_control='1') else v_message(1271 downto 1268);
   v_message_align(1347 downto 1344)<=ch_message_align(1287 downto 1284) when (mux_control='1') else v_message(1287 downto 1284);
   v_message_align(1351 downto 1348)<=ch_message_align(1303 downto 1300) when (mux_control='1') else v_message(1303 downto 1300);
   v_message_align(1355 downto 1352)<=ch_message_align(1319 downto 1316) when (mux_control='1') else v_message(1319 downto 1316);
   v_message_align(1359 downto 1356)<=ch_message_align(1335 downto 1332) when (mux_control='1') else v_message(1335 downto 1332);
   v_message_align(1363 downto 1360)<=ch_message_align(1351 downto 1348) when (mux_control='1') else v_message(1351 downto 1348);
   v_message_align(1367 downto 1364)<=ch_message_align(1367 downto 1364) when (mux_control='1') else v_message(1367 downto 1364);
   v_message_align(1371 downto 1368)<=ch_message_align(1383 downto 1380) when (mux_control='1') else v_message(1383 downto 1380);
   v_message_align(1375 downto 1372)<=ch_message_align(1399 downto 1396) when (mux_control='1') else v_message(1399 downto 1396);
   v_message_align(1379 downto 1376)<=ch_message_align(1415 downto 1412) when (mux_control='1') else v_message(1415 downto 1412);
   v_message_align(1383 downto 1380)<=ch_message_align(1431 downto 1428) when (mux_control='1') else v_message(1431 downto 1428);
   v_message_align(1387 downto 1384)<=ch_message_align(1447 downto 1444) when (mux_control='1') else v_message(1447 downto 1444);
   v_message_align(1391 downto 1388)<=ch_message_align(1463 downto 1460) when (mux_control='1') else v_message(1463 downto 1460);
   v_message_align(1395 downto 1392)<=ch_message_align(1479 downto 1476) when (mux_control='1') else v_message(1479 downto 1476);
   v_message_align(1399 downto 1396)<=ch_message_align(1495 downto 1492) when (mux_control='1') else v_message(1495 downto 1492);
   v_message_align(1403 downto 1400)<=ch_message_align(1511 downto 1508) when (mux_control='1') else v_message(1511 downto 1508);
   v_message_align(1407 downto 1404)<=ch_message_align(1527 downto 1524) when (mux_control='1') else v_message(1527 downto 1524);
   v_message_align(1411 downto 1408)<=ch_message_align(1543 downto 1540) when (mux_control='1') else v_message(1543 downto 1540);
   v_message_align(1415 downto 1412)<=ch_message_align(1559 downto 1556) when (mux_control='1') else v_message(1559 downto 1556);
   v_message_align(1419 downto 1416)<=ch_message_align(1575 downto 1572) when (mux_control='1') else v_message(1575 downto 1572);
   v_message_align(1423 downto 1420)<=ch_message_align(1591 downto 1588) when (mux_control='1') else v_message(1591 downto 1588);
   v_message_align(1427 downto 1424)<=ch_message_align(1607 downto 1604) when (mux_control='1') else v_message(1607 downto 1604);
   v_message_align(1431 downto 1428)<=ch_message_align(1623 downto 1620) when (mux_control='1') else v_message(1623 downto 1620);
   v_message_align(1435 downto 1432)<=ch_message_align(1639 downto 1636) when (mux_control='1') else v_message(1639 downto 1636);
   v_message_align(1439 downto 1436)<=ch_message_align(1655 downto 1652) when (mux_control='1') else v_message(1655 downto 1652);
   v_message_align(1443 downto 1440)<=ch_message_align(1671 downto 1668) when (mux_control='1') else v_message(1671 downto 1668);
   v_message_align(1447 downto 1444)<=ch_message_align(1687 downto 1684) when (mux_control='1') else v_message(1687 downto 1684);
   v_message_align(1451 downto 1448)<=ch_message_align(1703 downto 1700) when (mux_control='1') else v_message(1703 downto 1700);
   v_message_align(1455 downto 1452)<=ch_message_align(1719 downto 1716) when (mux_control='1') else v_message(1719 downto 1716);
   v_message_align(1459 downto 1456)<=ch_message_align(1735 downto 1732) when (mux_control='1') else v_message(1735 downto 1732);
   v_message_align(1463 downto 1460)<=ch_message_align(1751 downto 1748) when (mux_control='1') else v_message(1751 downto 1748);
   v_message_align(1467 downto 1464)<=ch_message_align(1767 downto 1764) when (mux_control='1') else v_message(1767 downto 1764);
   v_message_align(1471 downto 1468)<=ch_message_align(1783 downto 1780) when (mux_control='1') else v_message(1783 downto 1780);
   v_message_align(1475 downto 1472)<=ch_message_align(1799 downto 1796) when (mux_control='1') else v_message(1799 downto 1796);
   v_message_align(1479 downto 1476)<=ch_message_align(1815 downto 1812) when (mux_control='1') else v_message(1815 downto 1812);
   v_message_align(1483 downto 1480)<=ch_message_align(1831 downto 1828) when (mux_control='1') else v_message(1831 downto 1828);
   v_message_align(1487 downto 1484)<=ch_message_align(1847 downto 1844) when (mux_control='1') else v_message(1847 downto 1844);
   v_message_align(1491 downto 1488)<=ch_message_align(1863 downto 1860) when (mux_control='1') else v_message(1863 downto 1860);
   v_message_align(1495 downto 1492)<=ch_message_align(1879 downto 1876) when (mux_control='1') else v_message(1879 downto 1876);
   v_message_align(1499 downto 1496)<=ch_message_align(1895 downto 1892) when (mux_control='1') else v_message(1895 downto 1892);
   v_message_align(1503 downto 1500)<=ch_message_align(1911 downto 1908) when (mux_control='1') else v_message(1911 downto 1908);
   v_message_align(1507 downto 1504)<=ch_message_align(1927 downto 1924) when (mux_control='1') else v_message(1927 downto 1924);
   v_message_align(1511 downto 1508)<=ch_message_align(1943 downto 1940) when (mux_control='1') else v_message(1943 downto 1940);
   v_message_align(1515 downto 1512)<=ch_message_align(1959 downto 1956) when (mux_control='1') else v_message(1959 downto 1956);
   v_message_align(1519 downto 1516)<=ch_message_align(1975 downto 1972) when (mux_control='1') else v_message(1975 downto 1972);
   v_message_align(1523 downto 1520)<=ch_message_align(1991 downto 1988) when (mux_control='1') else v_message(1991 downto 1988);
   v_message_align(1527 downto 1524)<=ch_message_align(2007 downto 2004) when (mux_control='1') else v_message(2007 downto 2004);
   v_message_align(1531 downto 1528)<=ch_message_align(2023 downto 2020) when (mux_control='1') else v_message(2023 downto 2020);
   v_message_align(1535 downto 1532)<=ch_message_align(2039 downto 2036) when (mux_control='1') else v_message(2039 downto 2036);
   v_message_align(1539 downto 1536)<=ch_message_align(15 downto 12) when (mux_control='1') else v_message(15 downto 12);
   v_message_align(1543 downto 1540)<=ch_message_align(31 downto 28) when (mux_control='1') else v_message(31 downto 28);
   v_message_align(1547 downto 1544)<=ch_message_align(47 downto 44) when (mux_control='1') else v_message(47 downto 44);
   v_message_align(1551 downto 1548)<=ch_message_align(63 downto 60) when (mux_control='1') else v_message(63 downto 60);
   v_message_align(1555 downto 1552)<=ch_message_align(79 downto 76) when (mux_control='1') else v_message(79 downto 76);
   v_message_align(1559 downto 1556)<=ch_message_align(95 downto 92) when (mux_control='1') else v_message(95 downto 92);
   v_message_align(1563 downto 1560)<=ch_message_align(111 downto 108) when (mux_control='1') else v_message(111 downto 108);
   v_message_align(1567 downto 1564)<=ch_message_align(127 downto 124) when (mux_control='1') else v_message(127 downto 124);
   v_message_align(1571 downto 1568)<=ch_message_align(143 downto 140) when (mux_control='1') else v_message(143 downto 140);
   v_message_align(1575 downto 1572)<=ch_message_align(159 downto 156) when (mux_control='1') else v_message(159 downto 156);
   v_message_align(1579 downto 1576)<=ch_message_align(175 downto 172) when (mux_control='1') else v_message(175 downto 172);
   v_message_align(1583 downto 1580)<=ch_message_align(191 downto 188) when (mux_control='1') else v_message(191 downto 188);
   v_message_align(1587 downto 1584)<=ch_message_align(207 downto 204) when (mux_control='1') else v_message(207 downto 204);
   v_message_align(1591 downto 1588)<=ch_message_align(223 downto 220) when (mux_control='1') else v_message(223 downto 220);
   v_message_align(1595 downto 1592)<=ch_message_align(239 downto 236) when (mux_control='1') else v_message(239 downto 236);
   v_message_align(1599 downto 1596)<=ch_message_align(255 downto 252) when (mux_control='1') else v_message(255 downto 252);
   v_message_align(1603 downto 1600)<=ch_message_align(271 downto 268) when (mux_control='1') else v_message(271 downto 268);
   v_message_align(1607 downto 1604)<=ch_message_align(287 downto 284) when (mux_control='1') else v_message(287 downto 284);
   v_message_align(1611 downto 1608)<=ch_message_align(303 downto 300) when (mux_control='1') else v_message(303 downto 300);
   v_message_align(1615 downto 1612)<=ch_message_align(319 downto 316) when (mux_control='1') else v_message(319 downto 316);
   v_message_align(1619 downto 1616)<=ch_message_align(335 downto 332) when (mux_control='1') else v_message(335 downto 332);
   v_message_align(1623 downto 1620)<=ch_message_align(351 downto 348) when (mux_control='1') else v_message(351 downto 348);
   v_message_align(1627 downto 1624)<=ch_message_align(367 downto 364) when (mux_control='1') else v_message(367 downto 364);
   v_message_align(1631 downto 1628)<=ch_message_align(383 downto 380) when (mux_control='1') else v_message(383 downto 380);
   v_message_align(1635 downto 1632)<=ch_message_align(399 downto 396) when (mux_control='1') else v_message(399 downto 396);
   v_message_align(1639 downto 1636)<=ch_message_align(415 downto 412) when (mux_control='1') else v_message(415 downto 412);
   v_message_align(1643 downto 1640)<=ch_message_align(431 downto 428) when (mux_control='1') else v_message(431 downto 428);
   v_message_align(1647 downto 1644)<=ch_message_align(447 downto 444) when (mux_control='1') else v_message(447 downto 444);
   v_message_align(1651 downto 1648)<=ch_message_align(463 downto 460) when (mux_control='1') else v_message(463 downto 460);
   v_message_align(1655 downto 1652)<=ch_message_align(479 downto 476) when (mux_control='1') else v_message(479 downto 476);
   v_message_align(1659 downto 1656)<=ch_message_align(495 downto 492) when (mux_control='1') else v_message(495 downto 492);
   v_message_align(1663 downto 1660)<=ch_message_align(511 downto 508) when (mux_control='1') else v_message(511 downto 508);
   v_message_align(1667 downto 1664)<=ch_message_align(527 downto 524) when (mux_control='1') else v_message(527 downto 524);
   v_message_align(1671 downto 1668)<=ch_message_align(543 downto 540) when (mux_control='1') else v_message(543 downto 540);
   v_message_align(1675 downto 1672)<=ch_message_align(559 downto 556) when (mux_control='1') else v_message(559 downto 556);
   v_message_align(1679 downto 1676)<=ch_message_align(575 downto 572) when (mux_control='1') else v_message(575 downto 572);
   v_message_align(1683 downto 1680)<=ch_message_align(591 downto 588) when (mux_control='1') else v_message(591 downto 588);
   v_message_align(1687 downto 1684)<=ch_message_align(607 downto 604) when (mux_control='1') else v_message(607 downto 604);
   v_message_align(1691 downto 1688)<=ch_message_align(623 downto 620) when (mux_control='1') else v_message(623 downto 620);
   v_message_align(1695 downto 1692)<=ch_message_align(639 downto 636) when (mux_control='1') else v_message(639 downto 636);
   v_message_align(1699 downto 1696)<=ch_message_align(655 downto 652) when (mux_control='1') else v_message(655 downto 652);
   v_message_align(1703 downto 1700)<=ch_message_align(671 downto 668) when (mux_control='1') else v_message(671 downto 668);
   v_message_align(1707 downto 1704)<=ch_message_align(687 downto 684) when (mux_control='1') else v_message(687 downto 684);
   v_message_align(1711 downto 1708)<=ch_message_align(703 downto 700) when (mux_control='1') else v_message(703 downto 700);
   v_message_align(1715 downto 1712)<=ch_message_align(719 downto 716) when (mux_control='1') else v_message(719 downto 716);
   v_message_align(1719 downto 1716)<=ch_message_align(735 downto 732) when (mux_control='1') else v_message(735 downto 732);
   v_message_align(1723 downto 1720)<=ch_message_align(751 downto 748) when (mux_control='1') else v_message(751 downto 748);
   v_message_align(1727 downto 1724)<=ch_message_align(767 downto 764) when (mux_control='1') else v_message(767 downto 764);
   v_message_align(1731 downto 1728)<=ch_message_align(783 downto 780) when (mux_control='1') else v_message(783 downto 780);
   v_message_align(1735 downto 1732)<=ch_message_align(799 downto 796) when (mux_control='1') else v_message(799 downto 796);
   v_message_align(1739 downto 1736)<=ch_message_align(815 downto 812) when (mux_control='1') else v_message(815 downto 812);
   v_message_align(1743 downto 1740)<=ch_message_align(831 downto 828) when (mux_control='1') else v_message(831 downto 828);
   v_message_align(1747 downto 1744)<=ch_message_align(847 downto 844) when (mux_control='1') else v_message(847 downto 844);
   v_message_align(1751 downto 1748)<=ch_message_align(863 downto 860) when (mux_control='1') else v_message(863 downto 860);
   v_message_align(1755 downto 1752)<=ch_message_align(879 downto 876) when (mux_control='1') else v_message(879 downto 876);
   v_message_align(1759 downto 1756)<=ch_message_align(895 downto 892) when (mux_control='1') else v_message(895 downto 892);
   v_message_align(1763 downto 1760)<=ch_message_align(911 downto 908) when (mux_control='1') else v_message(911 downto 908);
   v_message_align(1767 downto 1764)<=ch_message_align(927 downto 924) when (mux_control='1') else v_message(927 downto 924);
   v_message_align(1771 downto 1768)<=ch_message_align(943 downto 940) when (mux_control='1') else v_message(943 downto 940);
   v_message_align(1775 downto 1772)<=ch_message_align(959 downto 956) when (mux_control='1') else v_message(959 downto 956);
   v_message_align(1779 downto 1776)<=ch_message_align(975 downto 972) when (mux_control='1') else v_message(975 downto 972);
   v_message_align(1783 downto 1780)<=ch_message_align(991 downto 988) when (mux_control='1') else v_message(991 downto 988);
   v_message_align(1787 downto 1784)<=ch_message_align(1007 downto 1004) when (mux_control='1') else v_message(1007 downto 1004);
   v_message_align(1791 downto 1788)<=ch_message_align(1023 downto 1020) when (mux_control='1') else v_message(1023 downto 1020);
   v_message_align(1795 downto 1792)<=ch_message_align(1039 downto 1036) when (mux_control='1') else v_message(1039 downto 1036);
   v_message_align(1799 downto 1796)<=ch_message_align(1055 downto 1052) when (mux_control='1') else v_message(1055 downto 1052);
   v_message_align(1803 downto 1800)<=ch_message_align(1071 downto 1068) when (mux_control='1') else v_message(1071 downto 1068);
   v_message_align(1807 downto 1804)<=ch_message_align(1087 downto 1084) when (mux_control='1') else v_message(1087 downto 1084);
   v_message_align(1811 downto 1808)<=ch_message_align(1103 downto 1100) when (mux_control='1') else v_message(1103 downto 1100);
   v_message_align(1815 downto 1812)<=ch_message_align(1119 downto 1116) when (mux_control='1') else v_message(1119 downto 1116);
   v_message_align(1819 downto 1816)<=ch_message_align(1135 downto 1132) when (mux_control='1') else v_message(1135 downto 1132);
   v_message_align(1823 downto 1820)<=ch_message_align(1151 downto 1148) when (mux_control='1') else v_message(1151 downto 1148);
   v_message_align(1827 downto 1824)<=ch_message_align(1167 downto 1164) when (mux_control='1') else v_message(1167 downto 1164);
   v_message_align(1831 downto 1828)<=ch_message_align(1183 downto 1180) when (mux_control='1') else v_message(1183 downto 1180);
   v_message_align(1835 downto 1832)<=ch_message_align(1199 downto 1196) when (mux_control='1') else v_message(1199 downto 1196);
   v_message_align(1839 downto 1836)<=ch_message_align(1215 downto 1212) when (mux_control='1') else v_message(1215 downto 1212);
   v_message_align(1843 downto 1840)<=ch_message_align(1231 downto 1228) when (mux_control='1') else v_message(1231 downto 1228);
   v_message_align(1847 downto 1844)<=ch_message_align(1247 downto 1244) when (mux_control='1') else v_message(1247 downto 1244);
   v_message_align(1851 downto 1848)<=ch_message_align(1263 downto 1260) when (mux_control='1') else v_message(1263 downto 1260);
   v_message_align(1855 downto 1852)<=ch_message_align(1279 downto 1276) when (mux_control='1') else v_message(1279 downto 1276);
   v_message_align(1859 downto 1856)<=ch_message_align(1295 downto 1292) when (mux_control='1') else v_message(1295 downto 1292);
   v_message_align(1863 downto 1860)<=ch_message_align(1311 downto 1308) when (mux_control='1') else v_message(1311 downto 1308);
   v_message_align(1867 downto 1864)<=ch_message_align(1327 downto 1324) when (mux_control='1') else v_message(1327 downto 1324);
   v_message_align(1871 downto 1868)<=ch_message_align(1343 downto 1340) when (mux_control='1') else v_message(1343 downto 1340);
   v_message_align(1875 downto 1872)<=ch_message_align(1359 downto 1356) when (mux_control='1') else v_message(1359 downto 1356);
   v_message_align(1879 downto 1876)<=ch_message_align(1375 downto 1372) when (mux_control='1') else v_message(1375 downto 1372);
   v_message_align(1883 downto 1880)<=ch_message_align(1391 downto 1388) when (mux_control='1') else v_message(1391 downto 1388);
   v_message_align(1887 downto 1884)<=ch_message_align(1407 downto 1404) when (mux_control='1') else v_message(1407 downto 1404);
   v_message_align(1891 downto 1888)<=ch_message_align(1423 downto 1420) when (mux_control='1') else v_message(1423 downto 1420);
   v_message_align(1895 downto 1892)<=ch_message_align(1439 downto 1436) when (mux_control='1') else v_message(1439 downto 1436);
   v_message_align(1899 downto 1896)<=ch_message_align(1455 downto 1452) when (mux_control='1') else v_message(1455 downto 1452);
   v_message_align(1903 downto 1900)<=ch_message_align(1471 downto 1468) when (mux_control='1') else v_message(1471 downto 1468);
   v_message_align(1907 downto 1904)<=ch_message_align(1487 downto 1484) when (mux_control='1') else v_message(1487 downto 1484);
   v_message_align(1911 downto 1908)<=ch_message_align(1503 downto 1500) when (mux_control='1') else v_message(1503 downto 1500);
   v_message_align(1915 downto 1912)<=ch_message_align(1519 downto 1516) when (mux_control='1') else v_message(1519 downto 1516);
   v_message_align(1919 downto 1916)<=ch_message_align(1535 downto 1532) when (mux_control='1') else v_message(1535 downto 1532);
   v_message_align(1923 downto 1920)<=ch_message_align(1551 downto 1548) when (mux_control='1') else v_message(1551 downto 1548);
   v_message_align(1927 downto 1924)<=ch_message_align(1567 downto 1564) when (mux_control='1') else v_message(1567 downto 1564);
   v_message_align(1931 downto 1928)<=ch_message_align(1583 downto 1580) when (mux_control='1') else v_message(1583 downto 1580);
   v_message_align(1935 downto 1932)<=ch_message_align(1599 downto 1596) when (mux_control='1') else v_message(1599 downto 1596);
   v_message_align(1939 downto 1936)<=ch_message_align(1615 downto 1612) when (mux_control='1') else v_message(1615 downto 1612);
   v_message_align(1943 downto 1940)<=ch_message_align(1631 downto 1628) when (mux_control='1') else v_message(1631 downto 1628);
   v_message_align(1947 downto 1944)<=ch_message_align(1647 downto 1644) when (mux_control='1') else v_message(1647 downto 1644);
   v_message_align(1951 downto 1948)<=ch_message_align(1663 downto 1660) when (mux_control='1') else v_message(1663 downto 1660);
   v_message_align(1955 downto 1952)<=ch_message_align(1679 downto 1676) when (mux_control='1') else v_message(1679 downto 1676);
   v_message_align(1959 downto 1956)<=ch_message_align(1695 downto 1692) when (mux_control='1') else v_message(1695 downto 1692);
   v_message_align(1963 downto 1960)<=ch_message_align(1711 downto 1708) when (mux_control='1') else v_message(1711 downto 1708);
   v_message_align(1967 downto 1964)<=ch_message_align(1727 downto 1724) when (mux_control='1') else v_message(1727 downto 1724);
   v_message_align(1971 downto 1968)<=ch_message_align(1743 downto 1740) when (mux_control='1') else v_message(1743 downto 1740);
   v_message_align(1975 downto 1972)<=ch_message_align(1759 downto 1756) when (mux_control='1') else v_message(1759 downto 1756);
   v_message_align(1979 downto 1976)<=ch_message_align(1775 downto 1772) when (mux_control='1') else v_message(1775 downto 1772);
   v_message_align(1983 downto 1980)<=ch_message_align(1791 downto 1788) when (mux_control='1') else v_message(1791 downto 1788);
   v_message_align(1987 downto 1984)<=ch_message_align(1807 downto 1804) when (mux_control='1') else v_message(1807 downto 1804);
   v_message_align(1991 downto 1988)<=ch_message_align(1823 downto 1820) when (mux_control='1') else v_message(1823 downto 1820);
   v_message_align(1995 downto 1992)<=ch_message_align(1839 downto 1836) when (mux_control='1') else v_message(1839 downto 1836);
   v_message_align(1999 downto 1996)<=ch_message_align(1855 downto 1852) when (mux_control='1') else v_message(1855 downto 1852);
   v_message_align(2003 downto 2000)<=ch_message_align(1871 downto 1868) when (mux_control='1') else v_message(1871 downto 1868);
   v_message_align(2007 downto 2004)<=ch_message_align(1887 downto 1884) when (mux_control='1') else v_message(1887 downto 1884);
   v_message_align(2011 downto 2008)<=ch_message_align(1903 downto 1900) when (mux_control='1') else v_message(1903 downto 1900);
   v_message_align(2015 downto 2012)<=ch_message_align(1919 downto 1916) when (mux_control='1') else v_message(1919 downto 1916);
   v_message_align(2019 downto 2016)<=ch_message_align(1935 downto 1932) when (mux_control='1') else v_message(1935 downto 1932);
   v_message_align(2023 downto 2020)<=ch_message_align(1951 downto 1948) when (mux_control='1') else v_message(1951 downto 1948);
   v_message_align(2027 downto 2024)<=ch_message_align(1967 downto 1964) when (mux_control='1') else v_message(1967 downto 1964);
   v_message_align(2031 downto 2028)<=ch_message_align(1983 downto 1980) when (mux_control='1') else v_message(1983 downto 1980);
   v_message_align(2035 downto 2032)<=ch_message_align(1999 downto 1996) when (mux_control='1') else v_message(1999 downto 1996);
   v_message_align(2039 downto 2036)<=ch_message_align(2015 downto 2012) when (mux_control='1') else v_message(2015 downto 2012);
   v_message_align(2043 downto 2040)<=ch_message_align(2031 downto 2028) when (mux_control='1') else v_message(2031 downto 2028);
   v_message_align(2047 downto 2044)<=ch_message_align(2047 downto 2044) when (mux_control='1') else v_message(2047 downto 2044);
  end rtl;