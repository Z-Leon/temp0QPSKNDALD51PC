library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity	c_message_walign	 is         
port(
	 c_message : in std_logic_vector(2047 downto 0);
	 c_message_align : out std_logic_vector(2047 downto 0)
	  );	 
end	c_message_walign;

architecture rtl of c_message_walign is
 begin
  c_message_align(3 downto 0) <= c_message(3 downto 0);
  c_message_align(7 downto 4) <= c_message(131 downto 128);
  c_message_align(11 downto 8) <= c_message(259 downto 256);
  c_message_align(15 downto 12) <= c_message(387 downto 384);
  c_message_align(19 downto 16) <= c_message(515 downto 512);
  c_message_align(23 downto 20) <= c_message(643 downto 640);
  c_message_align(27 downto 24) <= c_message(771 downto 768);
  c_message_align(31 downto 28) <= c_message(899 downto 896);
  c_message_align(35 downto 32) <= c_message(11 downto 8);
  c_message_align(39 downto 36) <= c_message(139 downto 136);
  c_message_align(43 downto 40) <= c_message(267 downto 264);
  c_message_align(47 downto 44) <= c_message(395 downto 392);
  c_message_align(51 downto 48) <= c_message(523 downto 520);
  c_message_align(55 downto 52) <= c_message(651 downto 648);
  c_message_align(59 downto 56) <= c_message(779 downto 776);
  c_message_align(63 downto 60) <= c_message(907 downto 904);
  c_message_align(67 downto 64) <= c_message(19 downto 16);
  c_message_align(71 downto 68) <= c_message(147 downto 144);
  c_message_align(75 downto 72) <= c_message(275 downto 272);
  c_message_align(79 downto 76) <= c_message(403 downto 400);
  c_message_align(83 downto 80) <= c_message(531 downto 528);
  c_message_align(87 downto 84) <= c_message(659 downto 656);
  c_message_align(91 downto 88) <= c_message(787 downto 784);
  c_message_align(95 downto 92) <= c_message(915 downto 912);
  c_message_align(99 downto 96) <= c_message(27 downto 24);
  c_message_align(103 downto 100) <= c_message(155 downto 152);
  c_message_align(107 downto 104) <= c_message(283 downto 280);
  c_message_align(111 downto 108) <= c_message(411 downto 408);
  c_message_align(115 downto 112) <= c_message(539 downto 536);
  c_message_align(119 downto 116) <= c_message(667 downto 664);
  c_message_align(123 downto 120) <= c_message(795 downto 792);
  c_message_align(127 downto 124) <= c_message(923 downto 920);
  c_message_align(131 downto 128) <= c_message(35 downto 32);
  c_message_align(135 downto 132) <= c_message(163 downto 160);
  c_message_align(139 downto 136) <= c_message(291 downto 288);
  c_message_align(143 downto 140) <= c_message(419 downto 416);
  c_message_align(147 downto 144) <= c_message(547 downto 544);
  c_message_align(151 downto 148) <= c_message(675 downto 672);
  c_message_align(155 downto 152) <= c_message(803 downto 800);
  c_message_align(159 downto 156) <= c_message(931 downto 928);
  c_message_align(163 downto 160) <= c_message(43 downto 40);
  c_message_align(167 downto 164) <= c_message(171 downto 168);
  c_message_align(171 downto 168) <= c_message(299 downto 296);
  c_message_align(175 downto 172) <= c_message(427 downto 424);
  c_message_align(179 downto 176) <= c_message(555 downto 552);
  c_message_align(183 downto 180) <= c_message(683 downto 680);
  c_message_align(187 downto 184) <= c_message(811 downto 808);
  c_message_align(191 downto 188) <= c_message(939 downto 936);
  c_message_align(195 downto 192) <= c_message(51 downto 48);
  c_message_align(199 downto 196) <= c_message(179 downto 176);
  c_message_align(203 downto 200) <= c_message(307 downto 304);
  c_message_align(207 downto 204) <= c_message(435 downto 432);
  c_message_align(211 downto 208) <= c_message(563 downto 560);
  c_message_align(215 downto 212) <= c_message(691 downto 688);
  c_message_align(219 downto 216) <= c_message(819 downto 816);
  c_message_align(223 downto 220) <= c_message(947 downto 944);
  c_message_align(227 downto 224) <= c_message(59 downto 56);
  c_message_align(231 downto 228) <= c_message(187 downto 184);
  c_message_align(235 downto 232) <= c_message(315 downto 312);
  c_message_align(239 downto 236) <= c_message(443 downto 440);
  c_message_align(243 downto 240) <= c_message(571 downto 568);
  c_message_align(247 downto 244) <= c_message(699 downto 696);
  c_message_align(251 downto 248) <= c_message(827 downto 824);
  c_message_align(255 downto 252) <= c_message(955 downto 952);
  c_message_align(259 downto 256) <= c_message(67 downto 64);
  c_message_align(263 downto 260) <= c_message(195 downto 192);
  c_message_align(267 downto 264) <= c_message(323 downto 320);
  c_message_align(271 downto 268) <= c_message(451 downto 448);
  c_message_align(275 downto 272) <= c_message(579 downto 576);
  c_message_align(279 downto 276) <= c_message(707 downto 704);
  c_message_align(283 downto 280) <= c_message(835 downto 832);
  c_message_align(287 downto 284) <= c_message(963 downto 960);
  c_message_align(291 downto 288) <= c_message(75 downto 72);
  c_message_align(295 downto 292) <= c_message(203 downto 200);
  c_message_align(299 downto 296) <= c_message(331 downto 328);
  c_message_align(303 downto 300) <= c_message(459 downto 456);
  c_message_align(307 downto 304) <= c_message(587 downto 584);
  c_message_align(311 downto 308) <= c_message(715 downto 712);
  c_message_align(315 downto 312) <= c_message(843 downto 840);
  c_message_align(319 downto 316) <= c_message(971 downto 968);
  c_message_align(323 downto 320) <= c_message(83 downto 80);
  c_message_align(327 downto 324) <= c_message(211 downto 208);
  c_message_align(331 downto 328) <= c_message(339 downto 336);
  c_message_align(335 downto 332) <= c_message(467 downto 464);
  c_message_align(339 downto 336) <= c_message(595 downto 592);
  c_message_align(343 downto 340) <= c_message(723 downto 720);
  c_message_align(347 downto 344) <= c_message(851 downto 848);
  c_message_align(351 downto 348) <= c_message(979 downto 976);
  c_message_align(355 downto 352) <= c_message(91 downto 88);
  c_message_align(359 downto 356) <= c_message(219 downto 216);
  c_message_align(363 downto 360) <= c_message(347 downto 344);
  c_message_align(367 downto 364) <= c_message(475 downto 472);
  c_message_align(371 downto 368) <= c_message(603 downto 600);
  c_message_align(375 downto 372) <= c_message(731 downto 728);
  c_message_align(379 downto 376) <= c_message(859 downto 856);
  c_message_align(383 downto 380) <= c_message(987 downto 984);
  c_message_align(387 downto 384) <= c_message(99 downto 96);
  c_message_align(391 downto 388) <= c_message(227 downto 224);
  c_message_align(395 downto 392) <= c_message(355 downto 352);
  c_message_align(399 downto 396) <= c_message(483 downto 480);
  c_message_align(403 downto 400) <= c_message(611 downto 608);
  c_message_align(407 downto 404) <= c_message(739 downto 736);
  c_message_align(411 downto 408) <= c_message(867 downto 864);
  c_message_align(415 downto 412) <= c_message(995 downto 992);
  c_message_align(419 downto 416) <= c_message(107 downto 104);
  c_message_align(423 downto 420) <= c_message(235 downto 232);
  c_message_align(427 downto 424) <= c_message(363 downto 360);
  c_message_align(431 downto 428) <= c_message(491 downto 488);
  c_message_align(435 downto 432) <= c_message(619 downto 616);
  c_message_align(439 downto 436) <= c_message(747 downto 744);
  c_message_align(443 downto 440) <= c_message(875 downto 872);
  c_message_align(447 downto 444) <= c_message(1003 downto 1000);
  c_message_align(451 downto 448) <= c_message(115 downto 112);
  c_message_align(455 downto 452) <= c_message(243 downto 240);
  c_message_align(459 downto 456) <= c_message(371 downto 368);
  c_message_align(463 downto 460) <= c_message(499 downto 496);
  c_message_align(467 downto 464) <= c_message(627 downto 624);
  c_message_align(471 downto 468) <= c_message(755 downto 752);
  c_message_align(475 downto 472) <= c_message(883 downto 880);
  c_message_align(479 downto 476) <= c_message(1011 downto 1008);
  c_message_align(483 downto 480) <= c_message(123 downto 120);
  c_message_align(487 downto 484) <= c_message(251 downto 248);
  c_message_align(491 downto 488) <= c_message(379 downto 376);
  c_message_align(495 downto 492) <= c_message(507 downto 504);
  c_message_align(499 downto 496) <= c_message(635 downto 632);
  c_message_align(503 downto 500) <= c_message(763 downto 760);
  c_message_align(507 downto 504) <= c_message(891 downto 888);
  c_message_align(511 downto 508) <= c_message(1019 downto 1016);
  c_message_align(515 downto 512) <= c_message(1027 downto 1024);
  c_message_align(519 downto 516) <= c_message(1155 downto 1152);
  c_message_align(523 downto 520) <= c_message(1283 downto 1280);
  c_message_align(527 downto 524) <= c_message(1411 downto 1408);
  c_message_align(531 downto 528) <= c_message(1539 downto 1536);
  c_message_align(535 downto 532) <= c_message(1667 downto 1664);
  c_message_align(539 downto 536) <= c_message(1795 downto 1792);
  c_message_align(543 downto 540) <= c_message(1923 downto 1920);
  c_message_align(547 downto 544) <= c_message(1035 downto 1032);
  c_message_align(551 downto 548) <= c_message(1163 downto 1160);
  c_message_align(555 downto 552) <= c_message(1291 downto 1288);
  c_message_align(559 downto 556) <= c_message(1419 downto 1416);
  c_message_align(563 downto 560) <= c_message(1547 downto 1544);
  c_message_align(567 downto 564) <= c_message(1675 downto 1672);
  c_message_align(571 downto 568) <= c_message(1803 downto 1800);
  c_message_align(575 downto 572) <= c_message(1931 downto 1928);
  c_message_align(579 downto 576) <= c_message(1043 downto 1040);
  c_message_align(583 downto 580) <= c_message(1171 downto 1168);
  c_message_align(587 downto 584) <= c_message(1299 downto 1296);
  c_message_align(591 downto 588) <= c_message(1427 downto 1424);
  c_message_align(595 downto 592) <= c_message(1555 downto 1552);
  c_message_align(599 downto 596) <= c_message(1683 downto 1680);
  c_message_align(603 downto 600) <= c_message(1811 downto 1808);
  c_message_align(607 downto 604) <= c_message(1939 downto 1936);
  c_message_align(611 downto 608) <= c_message(1051 downto 1048);
  c_message_align(615 downto 612) <= c_message(1179 downto 1176);
  c_message_align(619 downto 616) <= c_message(1307 downto 1304);
  c_message_align(623 downto 620) <= c_message(1435 downto 1432);
  c_message_align(627 downto 624) <= c_message(1563 downto 1560);
  c_message_align(631 downto 628) <= c_message(1691 downto 1688);
  c_message_align(635 downto 632) <= c_message(1819 downto 1816);
  c_message_align(639 downto 636) <= c_message(1947 downto 1944);
  c_message_align(643 downto 640) <= c_message(1059 downto 1056);
  c_message_align(647 downto 644) <= c_message(1187 downto 1184);
  c_message_align(651 downto 648) <= c_message(1315 downto 1312);
  c_message_align(655 downto 652) <= c_message(1443 downto 1440);
  c_message_align(659 downto 656) <= c_message(1571 downto 1568);
  c_message_align(663 downto 660) <= c_message(1699 downto 1696);
  c_message_align(667 downto 664) <= c_message(1827 downto 1824);
  c_message_align(671 downto 668) <= c_message(1955 downto 1952);
  c_message_align(675 downto 672) <= c_message(1067 downto 1064);
  c_message_align(679 downto 676) <= c_message(1195 downto 1192);
  c_message_align(683 downto 680) <= c_message(1323 downto 1320);
  c_message_align(687 downto 684) <= c_message(1451 downto 1448);
  c_message_align(691 downto 688) <= c_message(1579 downto 1576);
  c_message_align(695 downto 692) <= c_message(1707 downto 1704);
  c_message_align(699 downto 696) <= c_message(1835 downto 1832);
  c_message_align(703 downto 700) <= c_message(1963 downto 1960);
  c_message_align(707 downto 704) <= c_message(1075 downto 1072);
  c_message_align(711 downto 708) <= c_message(1203 downto 1200);
  c_message_align(715 downto 712) <= c_message(1331 downto 1328);
  c_message_align(719 downto 716) <= c_message(1459 downto 1456);
  c_message_align(723 downto 720) <= c_message(1587 downto 1584);
  c_message_align(727 downto 724) <= c_message(1715 downto 1712);
  c_message_align(731 downto 728) <= c_message(1843 downto 1840);
  c_message_align(735 downto 732) <= c_message(1971 downto 1968);
  c_message_align(739 downto 736) <= c_message(1083 downto 1080);
  c_message_align(743 downto 740) <= c_message(1211 downto 1208);
  c_message_align(747 downto 744) <= c_message(1339 downto 1336);
  c_message_align(751 downto 748) <= c_message(1467 downto 1464);
  c_message_align(755 downto 752) <= c_message(1595 downto 1592);
  c_message_align(759 downto 756) <= c_message(1723 downto 1720);
  c_message_align(763 downto 760) <= c_message(1851 downto 1848);
  c_message_align(767 downto 764) <= c_message(1979 downto 1976);
  c_message_align(771 downto 768) <= c_message(1091 downto 1088);
  c_message_align(775 downto 772) <= c_message(1219 downto 1216);
  c_message_align(779 downto 776) <= c_message(1347 downto 1344);
  c_message_align(783 downto 780) <= c_message(1475 downto 1472);
  c_message_align(787 downto 784) <= c_message(1603 downto 1600);
  c_message_align(791 downto 788) <= c_message(1731 downto 1728);
  c_message_align(795 downto 792) <= c_message(1859 downto 1856);
  c_message_align(799 downto 796) <= c_message(1987 downto 1984);
  c_message_align(803 downto 800) <= c_message(1099 downto 1096);
  c_message_align(807 downto 804) <= c_message(1227 downto 1224);
  c_message_align(811 downto 808) <= c_message(1355 downto 1352);
  c_message_align(815 downto 812) <= c_message(1483 downto 1480);
  c_message_align(819 downto 816) <= c_message(1611 downto 1608);
  c_message_align(823 downto 820) <= c_message(1739 downto 1736);
  c_message_align(827 downto 824) <= c_message(1867 downto 1864);
  c_message_align(831 downto 828) <= c_message(1995 downto 1992);
  c_message_align(835 downto 832) <= c_message(1107 downto 1104);
  c_message_align(839 downto 836) <= c_message(1235 downto 1232);
  c_message_align(843 downto 840) <= c_message(1363 downto 1360);
  c_message_align(847 downto 844) <= c_message(1491 downto 1488);
  c_message_align(851 downto 848) <= c_message(1619 downto 1616);
  c_message_align(855 downto 852) <= c_message(1747 downto 1744);
  c_message_align(859 downto 856) <= c_message(1875 downto 1872);
  c_message_align(863 downto 860) <= c_message(2003 downto 2000);
  c_message_align(867 downto 864) <= c_message(1115 downto 1112);
  c_message_align(871 downto 868) <= c_message(1243 downto 1240);
  c_message_align(875 downto 872) <= c_message(1371 downto 1368);
  c_message_align(879 downto 876) <= c_message(1499 downto 1496);
  c_message_align(883 downto 880) <= c_message(1627 downto 1624);
  c_message_align(887 downto 884) <= c_message(1755 downto 1752);
  c_message_align(891 downto 888) <= c_message(1883 downto 1880);
  c_message_align(895 downto 892) <= c_message(2011 downto 2008);
  c_message_align(899 downto 896) <= c_message(1123 downto 1120);
  c_message_align(903 downto 900) <= c_message(1251 downto 1248);
  c_message_align(907 downto 904) <= c_message(1379 downto 1376);
  c_message_align(911 downto 908) <= c_message(1507 downto 1504);
  c_message_align(915 downto 912) <= c_message(1635 downto 1632);
  c_message_align(919 downto 916) <= c_message(1763 downto 1760);
  c_message_align(923 downto 920) <= c_message(1891 downto 1888);
  c_message_align(927 downto 924) <= c_message(2019 downto 2016);
  c_message_align(931 downto 928) <= c_message(1131 downto 1128);
  c_message_align(935 downto 932) <= c_message(1259 downto 1256);
  c_message_align(939 downto 936) <= c_message(1387 downto 1384);
  c_message_align(943 downto 940) <= c_message(1515 downto 1512);
  c_message_align(947 downto 944) <= c_message(1643 downto 1640);
  c_message_align(951 downto 948) <= c_message(1771 downto 1768);
  c_message_align(955 downto 952) <= c_message(1899 downto 1896);
  c_message_align(959 downto 956) <= c_message(2027 downto 2024);
  c_message_align(963 downto 960) <= c_message(1139 downto 1136);
  c_message_align(967 downto 964) <= c_message(1267 downto 1264);
  c_message_align(971 downto 968) <= c_message(1395 downto 1392);
  c_message_align(975 downto 972) <= c_message(1523 downto 1520);
  c_message_align(979 downto 976) <= c_message(1651 downto 1648);
  c_message_align(983 downto 980) <= c_message(1779 downto 1776);
  c_message_align(987 downto 984) <= c_message(1907 downto 1904);
  c_message_align(991 downto 988) <= c_message(2035 downto 2032);
  c_message_align(995 downto 992) <= c_message(1147 downto 1144);
  c_message_align(999 downto 996) <= c_message(1275 downto 1272);
  c_message_align(1003 downto 1000) <= c_message(1403 downto 1400);
  c_message_align(1007 downto 1004) <= c_message(1531 downto 1528);
  c_message_align(1011 downto 1008) <= c_message(1659 downto 1656);
  c_message_align(1015 downto 1012) <= c_message(1787 downto 1784);
  c_message_align(1019 downto 1016) <= c_message(1915 downto 1912);
  c_message_align(1023 downto 1020) <= c_message(2043 downto 2040);
  c_message_align(1027 downto 1024) <= c_message(7 downto 4);
  c_message_align(1031 downto 1028) <= c_message(135 downto 132);
  c_message_align(1035 downto 1032) <= c_message(263 downto 260);
  c_message_align(1039 downto 1036) <= c_message(391 downto 388);
  c_message_align(1043 downto 1040) <= c_message(519 downto 516);
  c_message_align(1047 downto 1044) <= c_message(647 downto 644);
  c_message_align(1051 downto 1048) <= c_message(775 downto 772);
  c_message_align(1055 downto 1052) <= c_message(903 downto 900);
  c_message_align(1059 downto 1056) <= c_message(15 downto 12);
  c_message_align(1063 downto 1060) <= c_message(143 downto 140);
  c_message_align(1067 downto 1064) <= c_message(271 downto 268);
  c_message_align(1071 downto 1068) <= c_message(399 downto 396);
  c_message_align(1075 downto 1072) <= c_message(527 downto 524);
  c_message_align(1079 downto 1076) <= c_message(655 downto 652);
  c_message_align(1083 downto 1080) <= c_message(783 downto 780);
  c_message_align(1087 downto 1084) <= c_message(911 downto 908);
  c_message_align(1091 downto 1088) <= c_message(23 downto 20);
  c_message_align(1095 downto 1092) <= c_message(151 downto 148);
  c_message_align(1099 downto 1096) <= c_message(279 downto 276);
  c_message_align(1103 downto 1100) <= c_message(407 downto 404);
  c_message_align(1107 downto 1104) <= c_message(535 downto 532);
  c_message_align(1111 downto 1108) <= c_message(663 downto 660);
  c_message_align(1115 downto 1112) <= c_message(791 downto 788);
  c_message_align(1119 downto 1116) <= c_message(919 downto 916);
  c_message_align(1123 downto 1120) <= c_message(31 downto 28);
  c_message_align(1127 downto 1124) <= c_message(159 downto 156);
  c_message_align(1131 downto 1128) <= c_message(287 downto 284);
  c_message_align(1135 downto 1132) <= c_message(415 downto 412);
  c_message_align(1139 downto 1136) <= c_message(543 downto 540);
  c_message_align(1143 downto 1140) <= c_message(671 downto 668);
  c_message_align(1147 downto 1144) <= c_message(799 downto 796);
  c_message_align(1151 downto 1148) <= c_message(927 downto 924);
  c_message_align(1155 downto 1152) <= c_message(39 downto 36);
  c_message_align(1159 downto 1156) <= c_message(167 downto 164);
  c_message_align(1163 downto 1160) <= c_message(295 downto 292);
  c_message_align(1167 downto 1164) <= c_message(423 downto 420);
  c_message_align(1171 downto 1168) <= c_message(551 downto 548);
  c_message_align(1175 downto 1172) <= c_message(679 downto 676);
  c_message_align(1179 downto 1176) <= c_message(807 downto 804);
  c_message_align(1183 downto 1180) <= c_message(935 downto 932);
  c_message_align(1187 downto 1184) <= c_message(47 downto 44);
  c_message_align(1191 downto 1188) <= c_message(175 downto 172);
  c_message_align(1195 downto 1192) <= c_message(303 downto 300);
  c_message_align(1199 downto 1196) <= c_message(431 downto 428);
  c_message_align(1203 downto 1200) <= c_message(559 downto 556);
  c_message_align(1207 downto 1204) <= c_message(687 downto 684);
  c_message_align(1211 downto 1208) <= c_message(815 downto 812);
  c_message_align(1215 downto 1212) <= c_message(943 downto 940);
  c_message_align(1219 downto 1216) <= c_message(55 downto 52);
  c_message_align(1223 downto 1220) <= c_message(183 downto 180);
  c_message_align(1227 downto 1224) <= c_message(311 downto 308);
  c_message_align(1231 downto 1228) <= c_message(439 downto 436);
  c_message_align(1235 downto 1232) <= c_message(567 downto 564);
  c_message_align(1239 downto 1236) <= c_message(695 downto 692);
  c_message_align(1243 downto 1240) <= c_message(823 downto 820);
  c_message_align(1247 downto 1244) <= c_message(951 downto 948);
  c_message_align(1251 downto 1248) <= c_message(63 downto 60);
  c_message_align(1255 downto 1252) <= c_message(191 downto 188);
  c_message_align(1259 downto 1256) <= c_message(319 downto 316);
  c_message_align(1263 downto 1260) <= c_message(447 downto 444);
  c_message_align(1267 downto 1264) <= c_message(575 downto 572);
  c_message_align(1271 downto 1268) <= c_message(703 downto 700);
  c_message_align(1275 downto 1272) <= c_message(831 downto 828);
  c_message_align(1279 downto 1276) <= c_message(959 downto 956);
  c_message_align(1283 downto 1280) <= c_message(71 downto 68);
  c_message_align(1287 downto 1284) <= c_message(199 downto 196);
  c_message_align(1291 downto 1288) <= c_message(327 downto 324);
  c_message_align(1295 downto 1292) <= c_message(455 downto 452);
  c_message_align(1299 downto 1296) <= c_message(583 downto 580);
  c_message_align(1303 downto 1300) <= c_message(711 downto 708);
  c_message_align(1307 downto 1304) <= c_message(839 downto 836);
  c_message_align(1311 downto 1308) <= c_message(967 downto 964);
  c_message_align(1315 downto 1312) <= c_message(79 downto 76);
  c_message_align(1319 downto 1316) <= c_message(207 downto 204);
  c_message_align(1323 downto 1320) <= c_message(335 downto 332);
  c_message_align(1327 downto 1324) <= c_message(463 downto 460);
  c_message_align(1331 downto 1328) <= c_message(591 downto 588);
  c_message_align(1335 downto 1332) <= c_message(719 downto 716);
  c_message_align(1339 downto 1336) <= c_message(847 downto 844);
  c_message_align(1343 downto 1340) <= c_message(975 downto 972);
  c_message_align(1347 downto 1344) <= c_message(87 downto 84);
  c_message_align(1351 downto 1348) <= c_message(215 downto 212);
  c_message_align(1355 downto 1352) <= c_message(343 downto 340);
  c_message_align(1359 downto 1356) <= c_message(471 downto 468);
  c_message_align(1363 downto 1360) <= c_message(599 downto 596);
  c_message_align(1367 downto 1364) <= c_message(727 downto 724);
  c_message_align(1371 downto 1368) <= c_message(855 downto 852);
  c_message_align(1375 downto 1372) <= c_message(983 downto 980);
  c_message_align(1379 downto 1376) <= c_message(95 downto 92);
  c_message_align(1383 downto 1380) <= c_message(223 downto 220);
  c_message_align(1387 downto 1384) <= c_message(351 downto 348);
  c_message_align(1391 downto 1388) <= c_message(479 downto 476);
  c_message_align(1395 downto 1392) <= c_message(607 downto 604);
  c_message_align(1399 downto 1396) <= c_message(735 downto 732);
  c_message_align(1403 downto 1400) <= c_message(863 downto 860);
  c_message_align(1407 downto 1404) <= c_message(991 downto 988);
  c_message_align(1411 downto 1408) <= c_message(103 downto 100);
  c_message_align(1415 downto 1412) <= c_message(231 downto 228);
  c_message_align(1419 downto 1416) <= c_message(359 downto 356);
  c_message_align(1423 downto 1420) <= c_message(487 downto 484);
  c_message_align(1427 downto 1424) <= c_message(615 downto 612);
  c_message_align(1431 downto 1428) <= c_message(743 downto 740);
  c_message_align(1435 downto 1432) <= c_message(871 downto 868);
  c_message_align(1439 downto 1436) <= c_message(999 downto 996);
  c_message_align(1443 downto 1440) <= c_message(111 downto 108);
  c_message_align(1447 downto 1444) <= c_message(239 downto 236);
  c_message_align(1451 downto 1448) <= c_message(367 downto 364);
  c_message_align(1455 downto 1452) <= c_message(495 downto 492);
  c_message_align(1459 downto 1456) <= c_message(623 downto 620);
  c_message_align(1463 downto 1460) <= c_message(751 downto 748);
  c_message_align(1467 downto 1464) <= c_message(879 downto 876);
  c_message_align(1471 downto 1468) <= c_message(1007 downto 1004);
  c_message_align(1475 downto 1472) <= c_message(119 downto 116);
  c_message_align(1479 downto 1476) <= c_message(247 downto 244);
  c_message_align(1483 downto 1480) <= c_message(375 downto 372);
  c_message_align(1487 downto 1484) <= c_message(503 downto 500);
  c_message_align(1491 downto 1488) <= c_message(631 downto 628);
  c_message_align(1495 downto 1492) <= c_message(759 downto 756);
  c_message_align(1499 downto 1496) <= c_message(887 downto 884);
  c_message_align(1503 downto 1500) <= c_message(1015 downto 1012);
  c_message_align(1507 downto 1504) <= c_message(127 downto 124);
  c_message_align(1511 downto 1508) <= c_message(255 downto 252);
  c_message_align(1515 downto 1512) <= c_message(383 downto 380);
  c_message_align(1519 downto 1516) <= c_message(511 downto 508);
  c_message_align(1523 downto 1520) <= c_message(639 downto 636);
  c_message_align(1527 downto 1524) <= c_message(767 downto 764);
  c_message_align(1531 downto 1528) <= c_message(895 downto 892);
  c_message_align(1535 downto 1532) <= c_message(1023 downto 1020);
  c_message_align(1539 downto 1536) <= c_message(1031 downto 1028);
  c_message_align(1543 downto 1540) <= c_message(1159 downto 1156);
  c_message_align(1547 downto 1544) <= c_message(1287 downto 1284);
  c_message_align(1551 downto 1548) <= c_message(1415 downto 1412);
  c_message_align(1555 downto 1552) <= c_message(1543 downto 1540);
  c_message_align(1559 downto 1556) <= c_message(1671 downto 1668);
  c_message_align(1563 downto 1560) <= c_message(1799 downto 1796);
  c_message_align(1567 downto 1564) <= c_message(1927 downto 1924);
  c_message_align(1571 downto 1568) <= c_message(1039 downto 1036);
  c_message_align(1575 downto 1572) <= c_message(1167 downto 1164);
  c_message_align(1579 downto 1576) <= c_message(1295 downto 1292);
  c_message_align(1583 downto 1580) <= c_message(1423 downto 1420);
  c_message_align(1587 downto 1584) <= c_message(1551 downto 1548);
  c_message_align(1591 downto 1588) <= c_message(1679 downto 1676);
  c_message_align(1595 downto 1592) <= c_message(1807 downto 1804);
  c_message_align(1599 downto 1596) <= c_message(1935 downto 1932);
  c_message_align(1603 downto 1600) <= c_message(1047 downto 1044);
  c_message_align(1607 downto 1604) <= c_message(1175 downto 1172);
  c_message_align(1611 downto 1608) <= c_message(1303 downto 1300);
  c_message_align(1615 downto 1612) <= c_message(1431 downto 1428);
  c_message_align(1619 downto 1616) <= c_message(1559 downto 1556);
  c_message_align(1623 downto 1620) <= c_message(1687 downto 1684);
  c_message_align(1627 downto 1624) <= c_message(1815 downto 1812);
  c_message_align(1631 downto 1628) <= c_message(1943 downto 1940);
  c_message_align(1635 downto 1632) <= c_message(1055 downto 1052);
  c_message_align(1639 downto 1636) <= c_message(1183 downto 1180);
  c_message_align(1643 downto 1640) <= c_message(1311 downto 1308);
  c_message_align(1647 downto 1644) <= c_message(1439 downto 1436);
  c_message_align(1651 downto 1648) <= c_message(1567 downto 1564);
  c_message_align(1655 downto 1652) <= c_message(1695 downto 1692);
  c_message_align(1659 downto 1656) <= c_message(1823 downto 1820);
  c_message_align(1663 downto 1660) <= c_message(1951 downto 1948);
  c_message_align(1667 downto 1664) <= c_message(1063 downto 1060);
  c_message_align(1671 downto 1668) <= c_message(1191 downto 1188);
  c_message_align(1675 downto 1672) <= c_message(1319 downto 1316);
  c_message_align(1679 downto 1676) <= c_message(1447 downto 1444);
  c_message_align(1683 downto 1680) <= c_message(1575 downto 1572);
  c_message_align(1687 downto 1684) <= c_message(1703 downto 1700);
  c_message_align(1691 downto 1688) <= c_message(1831 downto 1828);
  c_message_align(1695 downto 1692) <= c_message(1959 downto 1956);
  c_message_align(1699 downto 1696) <= c_message(1071 downto 1068);
  c_message_align(1703 downto 1700) <= c_message(1199 downto 1196);
  c_message_align(1707 downto 1704) <= c_message(1327 downto 1324);
  c_message_align(1711 downto 1708) <= c_message(1455 downto 1452);
  c_message_align(1715 downto 1712) <= c_message(1583 downto 1580);
  c_message_align(1719 downto 1716) <= c_message(1711 downto 1708);
  c_message_align(1723 downto 1720) <= c_message(1839 downto 1836);
  c_message_align(1727 downto 1724) <= c_message(1967 downto 1964);
  c_message_align(1731 downto 1728) <= c_message(1079 downto 1076);
  c_message_align(1735 downto 1732) <= c_message(1207 downto 1204);
  c_message_align(1739 downto 1736) <= c_message(1335 downto 1332);
  c_message_align(1743 downto 1740) <= c_message(1463 downto 1460);
  c_message_align(1747 downto 1744) <= c_message(1591 downto 1588);
  c_message_align(1751 downto 1748) <= c_message(1719 downto 1716);
  c_message_align(1755 downto 1752) <= c_message(1847 downto 1844);
  c_message_align(1759 downto 1756) <= c_message(1975 downto 1972);
  c_message_align(1763 downto 1760) <= c_message(1087 downto 1084);
  c_message_align(1767 downto 1764) <= c_message(1215 downto 1212);
  c_message_align(1771 downto 1768) <= c_message(1343 downto 1340);
  c_message_align(1775 downto 1772) <= c_message(1471 downto 1468);
  c_message_align(1779 downto 1776) <= c_message(1599 downto 1596);
  c_message_align(1783 downto 1780) <= c_message(1727 downto 1724);
  c_message_align(1787 downto 1784) <= c_message(1855 downto 1852);
  c_message_align(1791 downto 1788) <= c_message(1983 downto 1980);
  c_message_align(1795 downto 1792) <= c_message(1095 downto 1092);
  c_message_align(1799 downto 1796) <= c_message(1223 downto 1220);
  c_message_align(1803 downto 1800) <= c_message(1351 downto 1348);
  c_message_align(1807 downto 1804) <= c_message(1479 downto 1476);
  c_message_align(1811 downto 1808) <= c_message(1607 downto 1604);
  c_message_align(1815 downto 1812) <= c_message(1735 downto 1732);
  c_message_align(1819 downto 1816) <= c_message(1863 downto 1860);
  c_message_align(1823 downto 1820) <= c_message(1991 downto 1988);
  c_message_align(1827 downto 1824) <= c_message(1103 downto 1100);
  c_message_align(1831 downto 1828) <= c_message(1231 downto 1228);
  c_message_align(1835 downto 1832) <= c_message(1359 downto 1356);
  c_message_align(1839 downto 1836) <= c_message(1487 downto 1484);
  c_message_align(1843 downto 1840) <= c_message(1615 downto 1612);
  c_message_align(1847 downto 1844) <= c_message(1743 downto 1740);
  c_message_align(1851 downto 1848) <= c_message(1871 downto 1868);
  c_message_align(1855 downto 1852) <= c_message(1999 downto 1996);
  c_message_align(1859 downto 1856) <= c_message(1111 downto 1108);
  c_message_align(1863 downto 1860) <= c_message(1239 downto 1236);
  c_message_align(1867 downto 1864) <= c_message(1367 downto 1364);
  c_message_align(1871 downto 1868) <= c_message(1495 downto 1492);
  c_message_align(1875 downto 1872) <= c_message(1623 downto 1620);
  c_message_align(1879 downto 1876) <= c_message(1751 downto 1748);
  c_message_align(1883 downto 1880) <= c_message(1879 downto 1876);
  c_message_align(1887 downto 1884) <= c_message(2007 downto 2004);
  c_message_align(1891 downto 1888) <= c_message(1119 downto 1116);
  c_message_align(1895 downto 1892) <= c_message(1247 downto 1244);
  c_message_align(1899 downto 1896) <= c_message(1375 downto 1372);
  c_message_align(1903 downto 1900) <= c_message(1503 downto 1500);
  c_message_align(1907 downto 1904) <= c_message(1631 downto 1628);
  c_message_align(1911 downto 1908) <= c_message(1759 downto 1756);
  c_message_align(1915 downto 1912) <= c_message(1887 downto 1884);
  c_message_align(1919 downto 1916) <= c_message(2015 downto 2012);
  c_message_align(1923 downto 1920) <= c_message(1127 downto 1124);
  c_message_align(1927 downto 1924) <= c_message(1255 downto 1252);
  c_message_align(1931 downto 1928) <= c_message(1383 downto 1380);
  c_message_align(1935 downto 1932) <= c_message(1511 downto 1508);
  c_message_align(1939 downto 1936) <= c_message(1639 downto 1636);
  c_message_align(1943 downto 1940) <= c_message(1767 downto 1764);
  c_message_align(1947 downto 1944) <= c_message(1895 downto 1892);
  c_message_align(1951 downto 1948) <= c_message(2023 downto 2020);
  c_message_align(1955 downto 1952) <= c_message(1135 downto 1132);
  c_message_align(1959 downto 1956) <= c_message(1263 downto 1260);
  c_message_align(1963 downto 1960) <= c_message(1391 downto 1388);
  c_message_align(1967 downto 1964) <= c_message(1519 downto 1516);
  c_message_align(1971 downto 1968) <= c_message(1647 downto 1644);
  c_message_align(1975 downto 1972) <= c_message(1775 downto 1772);
  c_message_align(1979 downto 1976) <= c_message(1903 downto 1900);
  c_message_align(1983 downto 1980) <= c_message(2031 downto 2028);
  c_message_align(1987 downto 1984) <= c_message(1143 downto 1140);
  c_message_align(1991 downto 1988) <= c_message(1271 downto 1268);
  c_message_align(1995 downto 1992) <= c_message(1399 downto 1396);
  c_message_align(1999 downto 1996) <= c_message(1527 downto 1524);
  c_message_align(2003 downto 2000) <= c_message(1655 downto 1652);
  c_message_align(2007 downto 2004) <= c_message(1783 downto 1780);
  c_message_align(2011 downto 2008) <= c_message(1911 downto 1908);
  c_message_align(2015 downto 2012) <= c_message(2039 downto 2036);
  c_message_align(2019 downto 2016) <= c_message(1151 downto 1148);
  c_message_align(2023 downto 2020) <= c_message(1279 downto 1276);
  c_message_align(2027 downto 2024) <= c_message(1407 downto 1404);
  c_message_align(2031 downto 2028) <= c_message(1535 downto 1532);
  c_message_align(2035 downto 2032) <= c_message(1663 downto 1660);
  c_message_align(2039 downto 2036) <= c_message(1791 downto 1788);
  c_message_align(2043 downto 2040) <= c_message(1919 downto 1916);
  c_message_align(2047 downto 2044) <= c_message(2047 downto 2044);  
 end rtl; 