LVDS_RX_32to64_inst : LVDS_RX_32to64 PORT MAP (
		rx_in	 => rx_in_sig,
		rx_inclock	 => rx_inclock_sig,
		rx_out	 => rx_out_sig
	);
