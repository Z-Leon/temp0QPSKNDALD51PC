--��������������������������������������������������������
--Author: Jiang Long (29-Sep-2014)
--����ʱ��Ƶ�ʱ����ϸ�Ϊ���ʱ��Ƶ�ʵ�1/3��
--�ϸ����������ת��ʱ��valid_out����ȷ
--��������������������������������������������������������
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity	P24toP8_14	is
	 generic(
		kDataWidth  : positive :=14 );
port(
		aReset	: in std_logic;
		clk_in		: in std_logic;
		clk_out		: in std_logic;
		data_in1		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in2		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in3		: in std_logic_vector(kDataWidth-1 downto 0);
		data_in4		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in5		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in6		: in std_logic_vector(kDataWidth-1 downto 0);
		data_in7		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in8		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in9		: in std_logic_vector(kDataWidth-1 downto 0);
		data_in10		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in11		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in12		: in std_logic_vector(kDataWidth-1 downto 0);
		data_in13		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in14		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in15		: in std_logic_vector(kDataWidth-1 downto 0);
		data_in16		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in17		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in18		: in std_logic_vector(kDataWidth-1 downto 0);
		data_in19		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in20		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in21		: in std_logic_vector(kDataWidth-1 downto 0);
		data_in22		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in23		: in std_logic_vector(kDataWidth-1 downto 0);
		--data_in24		: in std_logic_vector(kDataWidth-1 downto 0);
		--valid_in	: in std_logic;

		data_out1		: out std_logic_vector(kDataWidth-1 downto 0);
		data_out2		: out std_logic_vector(kDataWidth-1 downto 0);
		data_out3		: out std_logic_vector(kDataWidth-1 downto 0);
		data_out4		: out std_logic_vector(kDataWidth-1 downto 0);
		data_out5		: out std_logic_vector(kDataWidth-1 downto 0);
		data_out6		: out std_logic_vector(kDataWidth-1 downto 0);
		data_out7		: out std_logic_vector(kDataWidth-1 downto 0);
		data_out8		: out std_logic_vector(kDataWidth-1 downto 0)
		--valid_out	: out std_logic
		);
end	P24toP8_14;
architecture rtl of	P24toP8_14	is 
	type DataArray is array (natural range <>) of std_logic_vector(kDataWidth-1 downto 0);
	signal data_fifo: DataArray(71 downto 0);
	signal valid_fifo : std_logic_vector(71 downto 0);
	signal counter_in : integer range 0 to	2 := 0;
	signal counter_out : integer range 0 to	8 := 0;
begin
	--Process In
	process (aReset, clk_in)
	begin
		if aReset='1' then
			data_fifo(0)<=(others=>'0');
			--data_fifo(1)<=(others=>'0');
			--data_fifo(2)<=(others=>'0');
			data_fifo(3)<=(others=>'0');
			--data_fifo(4)<=(others=>'0');
			--data_fifo(5)<=(others=>'0');
			data_fifo(6)<=(others=>'0');
			--data_fifo(7)<=(others=>'0');
			--data_fifo(8)<=(others=>'0');
			data_fifo(9)<=(others=>'0');
			--data_fifo(10)<=(others=>'0');
			--data_fifo(11)<=(others=>'0');
			data_fifo(12)<=(others=>'0');
			--data_fifo(13)<=(others=>'0');
			--data_fifo(14)<=(others=>'0');
			data_fifo(15)<=(others=>'0');
			--data_fifo(16)<=(others=>'0');
			--data_fifo(17)<=(others=>'0');
			data_fifo(18)<=(others=>'0');
			--ata_fifo(19)<=(others=>'0');
			--data_fifo(20)<=(others=>'0');
			data_fifo(21)<=(others=>'0');
			--data_fifo(22)<=(others=>'0');
			--data_fifo(23)<=(others=>'0');
			data_fifo(24)<=(others=>'0');
			--ata_fifo(25)<=(others=>'0');
			--data_fifo(26)<=(others=>'0');
			data_fifo(27)<=(others=>'0');
			--data_fifo(28)<=(others=>'0');
			--data_fifo(29)<=(others=>'0');
			data_fifo(30)<=(others=>'0');
			--data_fifo(31)<=(others=>'0');
			--data_fifo(32)<=(others=>'0');
			data_fifo(33)<=(others=>'0');
			--data_fifo(34)<=(others=>'0');
			--data_fifo(35)<=(others=>'0');
			data_fifo(36)<=(others=>'0');
			--data_fifo(37)<=(others=>'0');
			--data_fifo(38)<=(others=>'0');
			data_fifo(39)<=(others=>'0');
			--data_fifo(40)<=(others=>'0');
			--data_fifo(41)<=(others=>'0');
			data_fifo(42)<=(others=>'0');
			--data_fifo(43)<=(others=>'0');
			--data_fifo(44)<=(others=>'0');
			data_fifo(45)<=(others=>'0');
			--data_fifo(46)<=(others=>'0');
			--data_fifo(47)<=(others=>'0');
			data_fifo(48)<=(others=>'0');
			--data_fifo(49)<=(others=>'0');
			--data_fifo(50)<=(others=>'0');
			data_fifo(51)<=(others=>'0');
			--data_fifo(52)<=(others=>'0');
			--data_fifo(53)<=(others=>'0');
			data_fifo(54)<=(others=>'0');
			--data_fifo(55)<=(others=>'0');
			--data_fifo(56)<=(others=>'0');
			data_fifo(57)<=(others=>'0');
			--data_fifo(58)<=(others=>'0');
			--data_fifo(59)<=(others=>'0');
			data_fifo(60)<=(others=>'0');
			--data_fifo(61)<=(others=>'0');
			--data_fifo(62)<=(others=>'0');
			data_fifo(63)<=(others=>'0');
			--data_fifo(64)<=(others=>'0');
			--data_fifo(65)<=(others=>'0');
			data_fifo(66)<=(others=>'0');
			--data_fifo(67)<=(others=>'0');
			--data_fifo(68)<=(others=>'0');
			data_fifo(69)<=(others=>'0');
			--data_fifo(70)<=(others=>'0');
			--data_fifo(71)<=(others=>'0');
			-- valid_fifo(0)<='0';
			-- valid_fifo(1)<='0';
			-- valid_fifo(2)<='0';
			-- valid_fifo(3)<='0';
			-- valid_fifo(4)<='0';
			-- valid_fifo(5)<='0';
			-- valid_fifo(6)<='0';
			-- valid_fifo(7)<='0';
			-- valid_fifo(8)<='0';
			-- valid_fifo(9)<='0';
			-- valid_fifo(10)<='0';
			-- valid_fifo(11)<='0';
			-- valid_fifo(12)<='0';
			-- valid_fifo(13)<='0';
			-- valid_fifo(14)<='0';
			-- valid_fifo(15)<='0';
			-- valid_fifo(16)<='0';
			-- valid_fifo(17)<='0';
			-- valid_fifo(18)<='0';
			-- valid_fifo(19)<='0';
			-- valid_fifo(20)<='0';
			-- valid_fifo(21)<='0';
			-- valid_fifo(22)<='0';
			-- valid_fifo(23)<='0';
			-- valid_fifo(24)<='0';
			-- valid_fifo(25)<='0';
			-- valid_fifo(26)<='0';
			-- valid_fifo(27)<='0';
			-- valid_fifo(28)<='0';
			-- valid_fifo(29)<='0';
			-- valid_fifo(30)<='0';
			-- valid_fifo(31)<='0';
			-- valid_fifo(32)<='0';
			-- valid_fifo(33)<='0';
			-- valid_fifo(34)<='0';
			-- valid_fifo(35)<='0';
			-- valid_fifo(36)<='0';
			-- valid_fifo(37)<='0';
			-- valid_fifo(38)<='0';
			-- valid_fifo(39)<='0';
			-- valid_fifo(40)<='0';
			-- valid_fifo(41)<='0';
			-- valid_fifo(42)<='0';
			-- valid_fifo(43)<='0';
			-- valid_fifo(44)<='0';
			-- valid_fifo(45)<='0';
			-- valid_fifo(46)<='0';
			-- valid_fifo(47)<='0';
			-- valid_fifo(48)<='0';
			-- valid_fifo(49)<='0';
			-- valid_fifo(50)<='0';
			-- valid_fifo(51)<='0';
			-- valid_fifo(52)<='0';
			-- valid_fifo(53)<='0';
			-- valid_fifo(54)<='0';
			-- valid_fifo(55)<='0';
			-- valid_fifo(56)<='0';
			-- valid_fifo(57)<='0';
			-- valid_fifo(58)<='0';
			-- valid_fifo(59)<='0';
			-- valid_fifo(60)<='0';
			-- valid_fifo(61)<='0';
			-- valid_fifo(62)<='0';
			-- valid_fifo(63)<='0';
			-- valid_fifo(64)<='0';
			-- valid_fifo(65)<='0';
			-- valid_fifo(66)<='0';
			-- valid_fifo(67)<='0';
			-- valid_fifo(68)<='0';
			-- valid_fifo(69)<='0';
			-- valid_fifo(70)<='0';
			-- valid_fifo(71)<='0';
			counter_in <= 0;
		elsif rising_edge(clk_in) then
			case counter_in is 
				when	0 =>
					data_fifo(24)<=data_in1;
					--data_fifo(25)<=data_in2;
					--data_fifo(26)<=data_in3;
					data_fifo(27)<=data_in4;
					--data_fifo(28)<=data_in5;
					--data_fifo(29)<=data_in6;
					data_fifo(30)<=data_in7;
					--data_fifo(31)<=data_in8;
					--data_fifo(32)<=data_in9;
					data_fifo(33)<=data_in10;
					--data_fifo(34)<=data_in11;
					--data_fifo(35)<=data_in12;
					data_fifo(36)<=data_in13;
					--data_fifo(37)<=data_in14;
					--data_fifo(38)<=data_in15;
					data_fifo(39)<=data_in16;
					--data_fifo(40)<=data_in17;
					--data_fifo(41)<=data_in18;
					data_fifo(42)<=data_in19;
					--data_fifo(43)<=data_in20;
					--data_fifo(44)<=data_in21;
					data_fifo(45)<=data_in22;
					--data_fifo(46)<=data_in23;
					--data_fifo(47)<=data_in24;
					-- valid_fifo(24)<=valid_in;
					-- valid_fifo(25)<=valid_in;
					-- valid_fifo(26)<=valid_in;
					-- valid_fifo(27)<=valid_in;
					-- valid_fifo(28)<=valid_in;
					-- valid_fifo(29)<=valid_in;
					-- valid_fifo(30)<=valid_in;
					-- valid_fifo(31)<=valid_in;
					-- valid_fifo(32)<=valid_in;
					-- valid_fifo(33)<=valid_in;
					-- valid_fifo(34)<=valid_in;
					-- valid_fifo(35)<=valid_in;
					-- valid_fifo(36)<=valid_in;
					-- valid_fifo(37)<=valid_in;
					-- valid_fifo(38)<=valid_in;
					-- valid_fifo(39)<=valid_in;
					-- valid_fifo(40)<=valid_in;
					-- valid_fifo(41)<=valid_in;
					-- valid_fifo(42)<=valid_in;
					-- valid_fifo(43)<=valid_in;
					-- valid_fifo(44)<=valid_in;
					-- valid_fifo(45)<=valid_in;
					-- valid_fifo(46)<=valid_in;
					-- valid_fifo(47)<=valid_in;
					counter_in<=1;
				when	1 =>
					data_fifo(48)<=data_in1;
					--data_fifo(49)<=data_in2;
					--data_fifo(50)<=data_in3;
					data_fifo(51)<=data_in4;
					--data_fifo(52)<=data_in5;
					--data_fifo(53)<=data_in6;
					data_fifo(54)<=data_in7;
					--data_fifo(55)<=data_in8;
					--data_fifo(56)<=data_in9;
					data_fifo(57)<=data_in10;
					--data_fifo(58)<=data_in11;
					--data_fifo(59)<=data_in12;
					data_fifo(60)<=data_in13;
					--data_fifo(61)<=data_in14;
					--data_fifo(62)<=data_in15;
					data_fifo(63)<=data_in16;
					--data_fifo(64)<=data_in17;
					--data_fifo(65)<=data_in18;
					data_fifo(66)<=data_in19;
					--data_fifo(67)<=data_in20;
					--data_fifo(68)<=data_in21;
					data_fifo(69)<=data_in22;
					--data_fifo(70)<=data_in23;
					--data_fifo(71)<=data_in24;
					-- valid_fifo(48)<=valid_in;
					-- valid_fifo(49)<=valid_in;
					-- valid_fifo(50)<=valid_in;
					-- valid_fifo(51)<=valid_in;
					-- valid_fifo(52)<=valid_in;
					-- valid_fifo(53)<=valid_in;
					-- valid_fifo(54)<=valid_in;
					-- valid_fifo(55)<=valid_in;
					-- valid_fifo(56)<=valid_in;
					-- valid_fifo(57)<=valid_in;
					-- valid_fifo(58)<=valid_in;
					-- valid_fifo(59)<=valid_in;
					-- valid_fifo(60)<=valid_in;
					-- valid_fifo(61)<=valid_in;
					-- valid_fifo(62)<=valid_in;
					-- valid_fifo(63)<=valid_in;
					-- valid_fifo(64)<=valid_in;
					-- valid_fifo(65)<=valid_in;
					-- valid_fifo(66)<=valid_in;
					-- valid_fifo(67)<=valid_in;
					-- valid_fifo(68)<=valid_in;
					-- valid_fifo(69)<=valid_in;
					-- valid_fifo(70)<=valid_in;
					-- valid_fifo(71)<=valid_in;
					counter_in<=2;
				when	2 =>
					data_fifo(0)<=data_in1;
					--data_fifo(1)<=data_in2;
					--data_fifo(2)<=data_in3;
					data_fifo(3)<=data_in4;
					--data_fifo(4)<=data_in5;
					--data_fifo(5)<=data_in6;
					data_fifo(6)<=data_in7;
					--data_fifo(7)<=data_in8;
					--data_fifo(8)<=data_in9;
					data_fifo(9)<=data_in10;
					--data_fifo(10)<=data_in11;
					--data_fifo(11)<=data_in12;
					data_fifo(12)<=data_in13;
					--data_fifo(13)<=data_in14;
					--data_fifo(14)<=data_in15;
					data_fifo(15)<=data_in16;
					--data_fifo(16)<=data_in17;
					--data_fifo(17)<=data_in18;
					data_fifo(18)<=data_in19;
					--data_fifo(19)<=data_in20;
					--data_fifo(20)<=data_in21;
					data_fifo(21)<=data_in22;
					--data_fifo(22)<=data_in23;
					--data_fifo(23)<=data_in24;
					-- valid_fifo(0)<=valid_in;
					-- valid_fifo(1)<=valid_in;
					-- valid_fifo(2)<=valid_in;
					-- valid_fifo(3)<=valid_in;
					-- valid_fifo(4)<=valid_in;
					-- valid_fifo(5)<=valid_in;
					-- valid_fifo(6)<=valid_in;
					-- valid_fifo(7)<=valid_in;
					-- valid_fifo(8)<=valid_in;
					-- valid_fifo(9)<=valid_in;
					-- valid_fifo(10)<=valid_in;
					-- valid_fifo(11)<=valid_in;
					-- valid_fifo(12)<=valid_in;
					-- valid_fifo(13)<=valid_in;
					-- valid_fifo(14)<=valid_in;
					-- valid_fifo(15)<=valid_in;
					-- valid_fifo(16)<=valid_in;
					-- valid_fifo(17)<=valid_in;
					-- valid_fifo(18)<=valid_in;
					-- valid_fifo(19)<=valid_in;
					-- valid_fifo(20)<=valid_in;
					-- valid_fifo(21)<=valid_in;
					-- valid_fifo(22)<=valid_in;
					-- valid_fifo(23)<=valid_in;
					counter_in<=0;
				when others =>
					null;
			end case;
		end if;
	end process;

	--Process Out
	process (aReset, clk_out)
	begin
		if aReset='1' then
			data_out1<=(others=>'0');
			data_out2<=(others=>'0');
			data_out3<=(others=>'0');
			data_out4<=(others=>'0');
			data_out5<=(others=>'0');
			data_out6<=(others=>'0');
			data_out7<=(others=>'0');
			data_out8<=(others=>'0');
			--valid_out<='0';
			counter_out <= 0;
		elsif rising_edge(clk_out) then
			case counter_out is 
				when	0 =>
					data_out1<=data_fifo(0);
					data_out2<=(others=>'0');
					data_out3<=(others=>'0');
					data_out4<=data_fifo(3);
					data_out5<=(others=>'0');
					data_out6<=(others=>'0');
					data_out7<=data_fifo(6);
					data_out8<=(others=>'0');
					--valid_out<=valid_fifo(0);
					counter_out<=1;
				when	1 =>
					data_out1<=(others=>'0');
					data_out2<=data_fifo(9);
					data_out3<=(others=>'0');
					data_out4<=(others=>'0');
					data_out5<=data_fifo(12);
					data_out6<=(others=>'0');
					data_out7<=(others=>'0');
					data_out8<=data_fifo(15);
					--valid_out<=valid_fifo(8);
					counter_out<=2;
				when	2 =>
					data_out1<=(others=>'0');
					data_out2<=(others=>'0');
					data_out3<=data_fifo(18);
					data_out4<=(others=>'0');
					data_out5<=(others=>'0');
					data_out6<=data_fifo(21);
					data_out7<=(others=>'0');
					data_out8<=(others=>'0');
					--valid_out<=valid_fifo(16);
					counter_out<=3;
				when	3 =>
					data_out1<=data_fifo(24);
					data_out2<=(others=>'0');
					data_out3<=(others=>'0');
					data_out4<=data_fifo(27);
					data_out5<=(others=>'0');
					data_out6<=(others=>'0');
					data_out7<=data_fifo(30);
					data_out8<=(others=>'0');
					--valid_out<=valid_fifo(24);
					counter_out<=4;
				when	4 =>
					data_out1<=(others=>'0');
					data_out2<=data_fifo(33);
					data_out3<=(others=>'0');
					data_out4<=(others=>'0');
					data_out5<=data_fifo(36);
					data_out6<=(others=>'0');
					data_out7<=(others=>'0');
					data_out8<=data_fifo(39);
					--valid_out<=valid_fifo(32);
					counter_out<=5;
				when	5 =>
					data_out1<=(others=>'0');
					data_out2<=(others=>'0');
					data_out3<=data_fifo(42);
					data_out4<=(others=>'0');
					data_out5<=(others=>'0');
					data_out6<=data_fifo(45);
					data_out7<=(others=>'0');
					data_out8<=(others=>'0');
					--valid_out<=valid_fifo(40);
					counter_out<=6;
				when	6 =>
					data_out1<=data_fifo(48);
					data_out2<=(others=>'0');
					data_out3<=(others=>'0');
					data_out4<=data_fifo(51);
					data_out5<=(others=>'0');
					data_out6<=(others=>'0');
					data_out7<=data_fifo(54);
					data_out8<=(others=>'0');
					--valid_out<=valid_fifo(48);
					counter_out<=7;
				when	7 =>
					data_out1<=(others=>'0');
					data_out2<=data_fifo(57);
					data_out3<=(others=>'0');
					data_out4<=(others=>'0');
					data_out5<=data_fifo(60);
					data_out6<=(others=>'0');
					data_out7<=(others=>'0');
					data_out8<=data_fifo(63);
					--valid_out<=valid_fifo(56);
					counter_out<=8;
				when	8 =>
					data_out1<=(others=>'0');
					data_out2<=(others=>'0');
					data_out3<=data_fifo(66);
					data_out4<=(others=>'0');
					data_out5<=(others=>'0');
					data_out6<=data_fifo(69);
					data_out7<=(others=>'0');
					data_out8<=(others=>'0');
					--valid_out<=valid_fifo(64);
					counter_out<=0;
				when others =>
					null;
			end case;
		end if;
	end process;
end rtl;
