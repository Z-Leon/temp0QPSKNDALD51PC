    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.std_logic_unsigned.all;
    use ieee.std_logic_arith.all;

	entity inforeg_7136 is
	port
	(
		reset     :  in std_logic;
		clk       :  in std_logic;
		
		info_in   :  in std_logic_vector(7 downto 0);
		info_val  :  in std_logic;
		info_ena  :  in std_logic;
		 
		inforeg   :  out std_logic_vector(7135 downto 0)
	);
	end inforeg_7136;
	
	architecture rtl of inforeg_7136 is
	
	signal temp_inforeg : std_logic_vector(7135 downto 0);

	begin
		inforeg <= temp_inforeg;
		
		process ( reset , clk )
		begin
			if ( reset = '1' ) then
				temp_inforeg <= (others=>'0');
			
			elsif rising_edge(clk) then
				if ((info_val = '1') and (info_ena = '1')) then
					temp_inforeg(7135 downto 7128) <= info_in;
					temp_inforeg(7127 downto 7120) <= temp_inforeg(7135 downto 7128);
					temp_inforeg(7119 downto 7112) <= temp_inforeg(7127 downto 7120);
					temp_inforeg(7111 downto 7104) <= temp_inforeg(7119 downto 7112);
					temp_inforeg(7103 downto 7096) <= temp_inforeg(7111 downto 7104);
					temp_inforeg(7095 downto 7088) <= temp_inforeg(7103 downto 7096);
					temp_inforeg(7087 downto 7080) <= temp_inforeg(7095 downto 7088);
					temp_inforeg(7079 downto 7072) <= temp_inforeg(7087 downto 7080);
					temp_inforeg(7071 downto 7064) <= temp_inforeg(7079 downto 7072);
					temp_inforeg(7063 downto 7056) <= temp_inforeg(7071 downto 7064);
					temp_inforeg(7055 downto 7048) <= temp_inforeg(7063 downto 7056);
					temp_inforeg(7047 downto 7040) <= temp_inforeg(7055 downto 7048);
					temp_inforeg(7039 downto 7032) <= temp_inforeg(7047 downto 7040);
					temp_inforeg(7031 downto 7024) <= temp_inforeg(7039 downto 7032);
					temp_inforeg(7023 downto 7016) <= temp_inforeg(7031 downto 7024);
					temp_inforeg(7015 downto 7008) <= temp_inforeg(7023 downto 7016);
					temp_inforeg(7007 downto 7000) <= temp_inforeg(7015 downto 7008);
					temp_inforeg(6999 downto 6992) <= temp_inforeg(7007 downto 7000);
					temp_inforeg(6991 downto 6984) <= temp_inforeg(6999 downto 6992);
					temp_inforeg(6983 downto 6976) <= temp_inforeg(6991 downto 6984);
					temp_inforeg(6975 downto 6968) <= temp_inforeg(6983 downto 6976);
					temp_inforeg(6967 downto 6960) <= temp_inforeg(6975 downto 6968);
					temp_inforeg(6959 downto 6952) <= temp_inforeg(6967 downto 6960);
					temp_inforeg(6951 downto 6944) <= temp_inforeg(6959 downto 6952);
					temp_inforeg(6943 downto 6936) <= temp_inforeg(6951 downto 6944);
					temp_inforeg(6935 downto 6928) <= temp_inforeg(6943 downto 6936);
					temp_inforeg(6927 downto 6920) <= temp_inforeg(6935 downto 6928);
					temp_inforeg(6919 downto 6912) <= temp_inforeg(6927 downto 6920);
					temp_inforeg(6911 downto 6904) <= temp_inforeg(6919 downto 6912);
					temp_inforeg(6903 downto 6896) <= temp_inforeg(6911 downto 6904);
					temp_inforeg(6895 downto 6888) <= temp_inforeg(6903 downto 6896);
					temp_inforeg(6887 downto 6880) <= temp_inforeg(6895 downto 6888);
					temp_inforeg(6879 downto 6872) <= temp_inforeg(6887 downto 6880);
					temp_inforeg(6871 downto 6864) <= temp_inforeg(6879 downto 6872);
					temp_inforeg(6863 downto 6856) <= temp_inforeg(6871 downto 6864);
					temp_inforeg(6855 downto 6848) <= temp_inforeg(6863 downto 6856);
					temp_inforeg(6847 downto 6840) <= temp_inforeg(6855 downto 6848);
					temp_inforeg(6839 downto 6832) <= temp_inforeg(6847 downto 6840);
					temp_inforeg(6831 downto 6824) <= temp_inforeg(6839 downto 6832);
					temp_inforeg(6823 downto 6816) <= temp_inforeg(6831 downto 6824);
					temp_inforeg(6815 downto 6808) <= temp_inforeg(6823 downto 6816);
					temp_inforeg(6807 downto 6800) <= temp_inforeg(6815 downto 6808);
					temp_inforeg(6799 downto 6792) <= temp_inforeg(6807 downto 6800);
					temp_inforeg(6791 downto 6784) <= temp_inforeg(6799 downto 6792);
					temp_inforeg(6783 downto 6776) <= temp_inforeg(6791 downto 6784);
					temp_inforeg(6775 downto 6768) <= temp_inforeg(6783 downto 6776);
					temp_inforeg(6767 downto 6760) <= temp_inforeg(6775 downto 6768);
					temp_inforeg(6759 downto 6752) <= temp_inforeg(6767 downto 6760);
					temp_inforeg(6751 downto 6744) <= temp_inforeg(6759 downto 6752);
					temp_inforeg(6743 downto 6736) <= temp_inforeg(6751 downto 6744);
					temp_inforeg(6735 downto 6728) <= temp_inforeg(6743 downto 6736);
					temp_inforeg(6727 downto 6720) <= temp_inforeg(6735 downto 6728);
					temp_inforeg(6719 downto 6712) <= temp_inforeg(6727 downto 6720);
					temp_inforeg(6711 downto 6704) <= temp_inforeg(6719 downto 6712);
					temp_inforeg(6703 downto 6696) <= temp_inforeg(6711 downto 6704);
					temp_inforeg(6695 downto 6688) <= temp_inforeg(6703 downto 6696);
					temp_inforeg(6687 downto 6680) <= temp_inforeg(6695 downto 6688);
					temp_inforeg(6679 downto 6672) <= temp_inforeg(6687 downto 6680);
					temp_inforeg(6671 downto 6664) <= temp_inforeg(6679 downto 6672);
					temp_inforeg(6663 downto 6656) <= temp_inforeg(6671 downto 6664);
					temp_inforeg(6655 downto 6648) <= temp_inforeg(6663 downto 6656);
					temp_inforeg(6647 downto 6640) <= temp_inforeg(6655 downto 6648);
					temp_inforeg(6639 downto 6632) <= temp_inforeg(6647 downto 6640);
					temp_inforeg(6631 downto 6624) <= temp_inforeg(6639 downto 6632);
					temp_inforeg(6623 downto 6616) <= temp_inforeg(6631 downto 6624);
					temp_inforeg(6615 downto 6608) <= temp_inforeg(6623 downto 6616);
					temp_inforeg(6607 downto 6600) <= temp_inforeg(6615 downto 6608);
					temp_inforeg(6599 downto 6592) <= temp_inforeg(6607 downto 6600);
					temp_inforeg(6591 downto 6584) <= temp_inforeg(6599 downto 6592);
					temp_inforeg(6583 downto 6576) <= temp_inforeg(6591 downto 6584);
					temp_inforeg(6575 downto 6568) <= temp_inforeg(6583 downto 6576);
					temp_inforeg(6567 downto 6560) <= temp_inforeg(6575 downto 6568);
					temp_inforeg(6559 downto 6552) <= temp_inforeg(6567 downto 6560);
					temp_inforeg(6551 downto 6544) <= temp_inforeg(6559 downto 6552);
					temp_inforeg(6543 downto 6536) <= temp_inforeg(6551 downto 6544);
					temp_inforeg(6535 downto 6528) <= temp_inforeg(6543 downto 6536);
					temp_inforeg(6527 downto 6520) <= temp_inforeg(6535 downto 6528);
					temp_inforeg(6519 downto 6512) <= temp_inforeg(6527 downto 6520);
					temp_inforeg(6511 downto 6504) <= temp_inforeg(6519 downto 6512);
					temp_inforeg(6503 downto 6496) <= temp_inforeg(6511 downto 6504);
					temp_inforeg(6495 downto 6488) <= temp_inforeg(6503 downto 6496);
					temp_inforeg(6487 downto 6480) <= temp_inforeg(6495 downto 6488);
					temp_inforeg(6479 downto 6472) <= temp_inforeg(6487 downto 6480);
					temp_inforeg(6471 downto 6464) <= temp_inforeg(6479 downto 6472);
					temp_inforeg(6463 downto 6456) <= temp_inforeg(6471 downto 6464);
					temp_inforeg(6455 downto 6448) <= temp_inforeg(6463 downto 6456);
					temp_inforeg(6447 downto 6440) <= temp_inforeg(6455 downto 6448);
					temp_inforeg(6439 downto 6432) <= temp_inforeg(6447 downto 6440);
					temp_inforeg(6431 downto 6424) <= temp_inforeg(6439 downto 6432);
					temp_inforeg(6423 downto 6416) <= temp_inforeg(6431 downto 6424);
					temp_inforeg(6415 downto 6408) <= temp_inforeg(6423 downto 6416);
					temp_inforeg(6407 downto 6400) <= temp_inforeg(6415 downto 6408);
					temp_inforeg(6399 downto 6392) <= temp_inforeg(6407 downto 6400);
					temp_inforeg(6391 downto 6384) <= temp_inforeg(6399 downto 6392);
					temp_inforeg(6383 downto 6376) <= temp_inforeg(6391 downto 6384);
					temp_inforeg(6375 downto 6368) <= temp_inforeg(6383 downto 6376);
					temp_inforeg(6367 downto 6360) <= temp_inforeg(6375 downto 6368);
					temp_inforeg(6359 downto 6352) <= temp_inforeg(6367 downto 6360);
					temp_inforeg(6351 downto 6344) <= temp_inforeg(6359 downto 6352);
					temp_inforeg(6343 downto 6336) <= temp_inforeg(6351 downto 6344);
					temp_inforeg(6335 downto 6328) <= temp_inforeg(6343 downto 6336);
					temp_inforeg(6327 downto 6320) <= temp_inforeg(6335 downto 6328);
					temp_inforeg(6319 downto 6312) <= temp_inforeg(6327 downto 6320);
					temp_inforeg(6311 downto 6304) <= temp_inforeg(6319 downto 6312);
					temp_inforeg(6303 downto 6296) <= temp_inforeg(6311 downto 6304);
					temp_inforeg(6295 downto 6288) <= temp_inforeg(6303 downto 6296);
					temp_inforeg(6287 downto 6280) <= temp_inforeg(6295 downto 6288);
					temp_inforeg(6279 downto 6272) <= temp_inforeg(6287 downto 6280);
					temp_inforeg(6271 downto 6264) <= temp_inforeg(6279 downto 6272);
					temp_inforeg(6263 downto 6256) <= temp_inforeg(6271 downto 6264);
					temp_inforeg(6255 downto 6248) <= temp_inforeg(6263 downto 6256);
					temp_inforeg(6247 downto 6240) <= temp_inforeg(6255 downto 6248);
					temp_inforeg(6239 downto 6232) <= temp_inforeg(6247 downto 6240);
					temp_inforeg(6231 downto 6224) <= temp_inforeg(6239 downto 6232);
					temp_inforeg(6223 downto 6216) <= temp_inforeg(6231 downto 6224);
					temp_inforeg(6215 downto 6208) <= temp_inforeg(6223 downto 6216);
					temp_inforeg(6207 downto 6200) <= temp_inforeg(6215 downto 6208);
					temp_inforeg(6199 downto 6192) <= temp_inforeg(6207 downto 6200);
					temp_inforeg(6191 downto 6184) <= temp_inforeg(6199 downto 6192);
					temp_inforeg(6183 downto 6176) <= temp_inforeg(6191 downto 6184);
					temp_inforeg(6175 downto 6168) <= temp_inforeg(6183 downto 6176);
					temp_inforeg(6167 downto 6160) <= temp_inforeg(6175 downto 6168);
					temp_inforeg(6159 downto 6152) <= temp_inforeg(6167 downto 6160);
					temp_inforeg(6151 downto 6144) <= temp_inforeg(6159 downto 6152);
					temp_inforeg(6143 downto 6136) <= temp_inforeg(6151 downto 6144);
					temp_inforeg(6135 downto 6128) <= temp_inforeg(6143 downto 6136);
					temp_inforeg(6127 downto 6120) <= temp_inforeg(6135 downto 6128);
					temp_inforeg(6119 downto 6112) <= temp_inforeg(6127 downto 6120);
					temp_inforeg(6111 downto 6104) <= temp_inforeg(6119 downto 6112);
					temp_inforeg(6103 downto 6096) <= temp_inforeg(6111 downto 6104);
					temp_inforeg(6095 downto 6088) <= temp_inforeg(6103 downto 6096);
					temp_inforeg(6087 downto 6080) <= temp_inforeg(6095 downto 6088);
					temp_inforeg(6079 downto 6072) <= temp_inforeg(6087 downto 6080);
					temp_inforeg(6071 downto 6064) <= temp_inforeg(6079 downto 6072);
					temp_inforeg(6063 downto 6056) <= temp_inforeg(6071 downto 6064);
					temp_inforeg(6055 downto 6048) <= temp_inforeg(6063 downto 6056);
					temp_inforeg(6047 downto 6040) <= temp_inforeg(6055 downto 6048);
					temp_inforeg(6039 downto 6032) <= temp_inforeg(6047 downto 6040);
					temp_inforeg(6031 downto 6024) <= temp_inforeg(6039 downto 6032);
					temp_inforeg(6023 downto 6016) <= temp_inforeg(6031 downto 6024);
					temp_inforeg(6015 downto 6008) <= temp_inforeg(6023 downto 6016);
					temp_inforeg(6007 downto 6000) <= temp_inforeg(6015 downto 6008);
					temp_inforeg(5999 downto 5992) <= temp_inforeg(6007 downto 6000);
					temp_inforeg(5991 downto 5984) <= temp_inforeg(5999 downto 5992);
					temp_inforeg(5983 downto 5976) <= temp_inforeg(5991 downto 5984);
					temp_inforeg(5975 downto 5968) <= temp_inforeg(5983 downto 5976);
					temp_inforeg(5967 downto 5960) <= temp_inforeg(5975 downto 5968);
					temp_inforeg(5959 downto 5952) <= temp_inforeg(5967 downto 5960);
					temp_inforeg(5951 downto 5944) <= temp_inforeg(5959 downto 5952);
					temp_inforeg(5943 downto 5936) <= temp_inforeg(5951 downto 5944);
					temp_inforeg(5935 downto 5928) <= temp_inforeg(5943 downto 5936);
					temp_inforeg(5927 downto 5920) <= temp_inforeg(5935 downto 5928);
					temp_inforeg(5919 downto 5912) <= temp_inforeg(5927 downto 5920);
					temp_inforeg(5911 downto 5904) <= temp_inforeg(5919 downto 5912);
					temp_inforeg(5903 downto 5896) <= temp_inforeg(5911 downto 5904);
					temp_inforeg(5895 downto 5888) <= temp_inforeg(5903 downto 5896);
					temp_inforeg(5887 downto 5880) <= temp_inforeg(5895 downto 5888);
					temp_inforeg(5879 downto 5872) <= temp_inforeg(5887 downto 5880);
					temp_inforeg(5871 downto 5864) <= temp_inforeg(5879 downto 5872);
					temp_inforeg(5863 downto 5856) <= temp_inforeg(5871 downto 5864);
					temp_inforeg(5855 downto 5848) <= temp_inforeg(5863 downto 5856);
					temp_inforeg(5847 downto 5840) <= temp_inforeg(5855 downto 5848);
					temp_inforeg(5839 downto 5832) <= temp_inforeg(5847 downto 5840);
					temp_inforeg(5831 downto 5824) <= temp_inforeg(5839 downto 5832);
					temp_inforeg(5823 downto 5816) <= temp_inforeg(5831 downto 5824);
					temp_inforeg(5815 downto 5808) <= temp_inforeg(5823 downto 5816);
					temp_inforeg(5807 downto 5800) <= temp_inforeg(5815 downto 5808);
					temp_inforeg(5799 downto 5792) <= temp_inforeg(5807 downto 5800);
					temp_inforeg(5791 downto 5784) <= temp_inforeg(5799 downto 5792);
					temp_inforeg(5783 downto 5776) <= temp_inforeg(5791 downto 5784);
					temp_inforeg(5775 downto 5768) <= temp_inforeg(5783 downto 5776);
					temp_inforeg(5767 downto 5760) <= temp_inforeg(5775 downto 5768);
					temp_inforeg(5759 downto 5752) <= temp_inforeg(5767 downto 5760);
					temp_inforeg(5751 downto 5744) <= temp_inforeg(5759 downto 5752);
					temp_inforeg(5743 downto 5736) <= temp_inforeg(5751 downto 5744);
					temp_inforeg(5735 downto 5728) <= temp_inforeg(5743 downto 5736);
					temp_inforeg(5727 downto 5720) <= temp_inforeg(5735 downto 5728);
					temp_inforeg(5719 downto 5712) <= temp_inforeg(5727 downto 5720);
					temp_inforeg(5711 downto 5704) <= temp_inforeg(5719 downto 5712);
					temp_inforeg(5703 downto 5696) <= temp_inforeg(5711 downto 5704);
					temp_inforeg(5695 downto 5688) <= temp_inforeg(5703 downto 5696);
					temp_inforeg(5687 downto 5680) <= temp_inforeg(5695 downto 5688);
					temp_inforeg(5679 downto 5672) <= temp_inforeg(5687 downto 5680);
					temp_inforeg(5671 downto 5664) <= temp_inforeg(5679 downto 5672);
					temp_inforeg(5663 downto 5656) <= temp_inforeg(5671 downto 5664);
					temp_inforeg(5655 downto 5648) <= temp_inforeg(5663 downto 5656);
					temp_inforeg(5647 downto 5640) <= temp_inforeg(5655 downto 5648);
					temp_inforeg(5639 downto 5632) <= temp_inforeg(5647 downto 5640);
					temp_inforeg(5631 downto 5624) <= temp_inforeg(5639 downto 5632);
					temp_inforeg(5623 downto 5616) <= temp_inforeg(5631 downto 5624);
					temp_inforeg(5615 downto 5608) <= temp_inforeg(5623 downto 5616);
					temp_inforeg(5607 downto 5600) <= temp_inforeg(5615 downto 5608);
					temp_inforeg(5599 downto 5592) <= temp_inforeg(5607 downto 5600);
					temp_inforeg(5591 downto 5584) <= temp_inforeg(5599 downto 5592);
					temp_inforeg(5583 downto 5576) <= temp_inforeg(5591 downto 5584);
					temp_inforeg(5575 downto 5568) <= temp_inforeg(5583 downto 5576);
					temp_inforeg(5567 downto 5560) <= temp_inforeg(5575 downto 5568);
					temp_inforeg(5559 downto 5552) <= temp_inforeg(5567 downto 5560);
					temp_inforeg(5551 downto 5544) <= temp_inforeg(5559 downto 5552);
					temp_inforeg(5543 downto 5536) <= temp_inforeg(5551 downto 5544);
					temp_inforeg(5535 downto 5528) <= temp_inforeg(5543 downto 5536);
					temp_inforeg(5527 downto 5520) <= temp_inforeg(5535 downto 5528);
					temp_inforeg(5519 downto 5512) <= temp_inforeg(5527 downto 5520);
					temp_inforeg(5511 downto 5504) <= temp_inforeg(5519 downto 5512);
					temp_inforeg(5503 downto 5496) <= temp_inforeg(5511 downto 5504);
					temp_inforeg(5495 downto 5488) <= temp_inforeg(5503 downto 5496);
					temp_inforeg(5487 downto 5480) <= temp_inforeg(5495 downto 5488);
					temp_inforeg(5479 downto 5472) <= temp_inforeg(5487 downto 5480);
					temp_inforeg(5471 downto 5464) <= temp_inforeg(5479 downto 5472);
					temp_inforeg(5463 downto 5456) <= temp_inforeg(5471 downto 5464);
					temp_inforeg(5455 downto 5448) <= temp_inforeg(5463 downto 5456);
					temp_inforeg(5447 downto 5440) <= temp_inforeg(5455 downto 5448);
					temp_inforeg(5439 downto 5432) <= temp_inforeg(5447 downto 5440);
					temp_inforeg(5431 downto 5424) <= temp_inforeg(5439 downto 5432);
					temp_inforeg(5423 downto 5416) <= temp_inforeg(5431 downto 5424);
					temp_inforeg(5415 downto 5408) <= temp_inforeg(5423 downto 5416);
					temp_inforeg(5407 downto 5400) <= temp_inforeg(5415 downto 5408);
					temp_inforeg(5399 downto 5392) <= temp_inforeg(5407 downto 5400);
					temp_inforeg(5391 downto 5384) <= temp_inforeg(5399 downto 5392);
					temp_inforeg(5383 downto 5376) <= temp_inforeg(5391 downto 5384);
					temp_inforeg(5375 downto 5368) <= temp_inforeg(5383 downto 5376);
					temp_inforeg(5367 downto 5360) <= temp_inforeg(5375 downto 5368);
					temp_inforeg(5359 downto 5352) <= temp_inforeg(5367 downto 5360);
					temp_inforeg(5351 downto 5344) <= temp_inforeg(5359 downto 5352);
					temp_inforeg(5343 downto 5336) <= temp_inforeg(5351 downto 5344);
					temp_inforeg(5335 downto 5328) <= temp_inforeg(5343 downto 5336);
					temp_inforeg(5327 downto 5320) <= temp_inforeg(5335 downto 5328);
					temp_inforeg(5319 downto 5312) <= temp_inforeg(5327 downto 5320);
					temp_inforeg(5311 downto 5304) <= temp_inforeg(5319 downto 5312);
					temp_inforeg(5303 downto 5296) <= temp_inforeg(5311 downto 5304);
					temp_inforeg(5295 downto 5288) <= temp_inforeg(5303 downto 5296);
					temp_inforeg(5287 downto 5280) <= temp_inforeg(5295 downto 5288);
					temp_inforeg(5279 downto 5272) <= temp_inforeg(5287 downto 5280);
					temp_inforeg(5271 downto 5264) <= temp_inforeg(5279 downto 5272);
					temp_inforeg(5263 downto 5256) <= temp_inforeg(5271 downto 5264);
					temp_inforeg(5255 downto 5248) <= temp_inforeg(5263 downto 5256);
					temp_inforeg(5247 downto 5240) <= temp_inforeg(5255 downto 5248);
					temp_inforeg(5239 downto 5232) <= temp_inforeg(5247 downto 5240);
					temp_inforeg(5231 downto 5224) <= temp_inforeg(5239 downto 5232);
					temp_inforeg(5223 downto 5216) <= temp_inforeg(5231 downto 5224);
					temp_inforeg(5215 downto 5208) <= temp_inforeg(5223 downto 5216);
					temp_inforeg(5207 downto 5200) <= temp_inforeg(5215 downto 5208);
					temp_inforeg(5199 downto 5192) <= temp_inforeg(5207 downto 5200);
					temp_inforeg(5191 downto 5184) <= temp_inforeg(5199 downto 5192);
					temp_inforeg(5183 downto 5176) <= temp_inforeg(5191 downto 5184);
					temp_inforeg(5175 downto 5168) <= temp_inforeg(5183 downto 5176);
					temp_inforeg(5167 downto 5160) <= temp_inforeg(5175 downto 5168);
					temp_inforeg(5159 downto 5152) <= temp_inforeg(5167 downto 5160);
					temp_inforeg(5151 downto 5144) <= temp_inforeg(5159 downto 5152);
					temp_inforeg(5143 downto 5136) <= temp_inforeg(5151 downto 5144);
					temp_inforeg(5135 downto 5128) <= temp_inforeg(5143 downto 5136);
					temp_inforeg(5127 downto 5120) <= temp_inforeg(5135 downto 5128);
					temp_inforeg(5119 downto 5112) <= temp_inforeg(5127 downto 5120);
					temp_inforeg(5111 downto 5104) <= temp_inforeg(5119 downto 5112);
					temp_inforeg(5103 downto 5096) <= temp_inforeg(5111 downto 5104);
					temp_inforeg(5095 downto 5088) <= temp_inforeg(5103 downto 5096);
					temp_inforeg(5087 downto 5080) <= temp_inforeg(5095 downto 5088);
					temp_inforeg(5079 downto 5072) <= temp_inforeg(5087 downto 5080);
					temp_inforeg(5071 downto 5064) <= temp_inforeg(5079 downto 5072);
					temp_inforeg(5063 downto 5056) <= temp_inforeg(5071 downto 5064);
					temp_inforeg(5055 downto 5048) <= temp_inforeg(5063 downto 5056);
					temp_inforeg(5047 downto 5040) <= temp_inforeg(5055 downto 5048);
					temp_inforeg(5039 downto 5032) <= temp_inforeg(5047 downto 5040);
					temp_inforeg(5031 downto 5024) <= temp_inforeg(5039 downto 5032);
					temp_inforeg(5023 downto 5016) <= temp_inforeg(5031 downto 5024);
					temp_inforeg(5015 downto 5008) <= temp_inforeg(5023 downto 5016);
					temp_inforeg(5007 downto 5000) <= temp_inforeg(5015 downto 5008);
					temp_inforeg(4999 downto 4992) <= temp_inforeg(5007 downto 5000);
					temp_inforeg(4991 downto 4984) <= temp_inforeg(4999 downto 4992);
					temp_inforeg(4983 downto 4976) <= temp_inforeg(4991 downto 4984);
					temp_inforeg(4975 downto 4968) <= temp_inforeg(4983 downto 4976);
					temp_inforeg(4967 downto 4960) <= temp_inforeg(4975 downto 4968);
					temp_inforeg(4959 downto 4952) <= temp_inforeg(4967 downto 4960);
					temp_inforeg(4951 downto 4944) <= temp_inforeg(4959 downto 4952);
					temp_inforeg(4943 downto 4936) <= temp_inforeg(4951 downto 4944);
					temp_inforeg(4935 downto 4928) <= temp_inforeg(4943 downto 4936);
					temp_inforeg(4927 downto 4920) <= temp_inforeg(4935 downto 4928);
					temp_inforeg(4919 downto 4912) <= temp_inforeg(4927 downto 4920);
					temp_inforeg(4911 downto 4904) <= temp_inforeg(4919 downto 4912);
					temp_inforeg(4903 downto 4896) <= temp_inforeg(4911 downto 4904);
					temp_inforeg(4895 downto 4888) <= temp_inforeg(4903 downto 4896);
					temp_inforeg(4887 downto 4880) <= temp_inforeg(4895 downto 4888);
					temp_inforeg(4879 downto 4872) <= temp_inforeg(4887 downto 4880);
					temp_inforeg(4871 downto 4864) <= temp_inforeg(4879 downto 4872);
					temp_inforeg(4863 downto 4856) <= temp_inforeg(4871 downto 4864);
					temp_inforeg(4855 downto 4848) <= temp_inforeg(4863 downto 4856);
					temp_inforeg(4847 downto 4840) <= temp_inforeg(4855 downto 4848);
					temp_inforeg(4839 downto 4832) <= temp_inforeg(4847 downto 4840);
					temp_inforeg(4831 downto 4824) <= temp_inforeg(4839 downto 4832);
					temp_inforeg(4823 downto 4816) <= temp_inforeg(4831 downto 4824);
					temp_inforeg(4815 downto 4808) <= temp_inforeg(4823 downto 4816);
					temp_inforeg(4807 downto 4800) <= temp_inforeg(4815 downto 4808);
					temp_inforeg(4799 downto 4792) <= temp_inforeg(4807 downto 4800);
					temp_inforeg(4791 downto 4784) <= temp_inforeg(4799 downto 4792);
					temp_inforeg(4783 downto 4776) <= temp_inforeg(4791 downto 4784);
					temp_inforeg(4775 downto 4768) <= temp_inforeg(4783 downto 4776);
					temp_inforeg(4767 downto 4760) <= temp_inforeg(4775 downto 4768);
					temp_inforeg(4759 downto 4752) <= temp_inforeg(4767 downto 4760);
					temp_inforeg(4751 downto 4744) <= temp_inforeg(4759 downto 4752);
					temp_inforeg(4743 downto 4736) <= temp_inforeg(4751 downto 4744);
					temp_inforeg(4735 downto 4728) <= temp_inforeg(4743 downto 4736);
					temp_inforeg(4727 downto 4720) <= temp_inforeg(4735 downto 4728);
					temp_inforeg(4719 downto 4712) <= temp_inforeg(4727 downto 4720);
					temp_inforeg(4711 downto 4704) <= temp_inforeg(4719 downto 4712);
					temp_inforeg(4703 downto 4696) <= temp_inforeg(4711 downto 4704);
					temp_inforeg(4695 downto 4688) <= temp_inforeg(4703 downto 4696);
					temp_inforeg(4687 downto 4680) <= temp_inforeg(4695 downto 4688);
					temp_inforeg(4679 downto 4672) <= temp_inforeg(4687 downto 4680);
					temp_inforeg(4671 downto 4664) <= temp_inforeg(4679 downto 4672);
					temp_inforeg(4663 downto 4656) <= temp_inforeg(4671 downto 4664);
					temp_inforeg(4655 downto 4648) <= temp_inforeg(4663 downto 4656);
					temp_inforeg(4647 downto 4640) <= temp_inforeg(4655 downto 4648);
					temp_inforeg(4639 downto 4632) <= temp_inforeg(4647 downto 4640);
					temp_inforeg(4631 downto 4624) <= temp_inforeg(4639 downto 4632);
					temp_inforeg(4623 downto 4616) <= temp_inforeg(4631 downto 4624);
					temp_inforeg(4615 downto 4608) <= temp_inforeg(4623 downto 4616);
					temp_inforeg(4607 downto 4600) <= temp_inforeg(4615 downto 4608);
					temp_inforeg(4599 downto 4592) <= temp_inforeg(4607 downto 4600);
					temp_inforeg(4591 downto 4584) <= temp_inforeg(4599 downto 4592);
					temp_inforeg(4583 downto 4576) <= temp_inforeg(4591 downto 4584);
					temp_inforeg(4575 downto 4568) <= temp_inforeg(4583 downto 4576);
					temp_inforeg(4567 downto 4560) <= temp_inforeg(4575 downto 4568);
					temp_inforeg(4559 downto 4552) <= temp_inforeg(4567 downto 4560);
					temp_inforeg(4551 downto 4544) <= temp_inforeg(4559 downto 4552);
					temp_inforeg(4543 downto 4536) <= temp_inforeg(4551 downto 4544);
					temp_inforeg(4535 downto 4528) <= temp_inforeg(4543 downto 4536);
					temp_inforeg(4527 downto 4520) <= temp_inforeg(4535 downto 4528);
					temp_inforeg(4519 downto 4512) <= temp_inforeg(4527 downto 4520);
					temp_inforeg(4511 downto 4504) <= temp_inforeg(4519 downto 4512);
					temp_inforeg(4503 downto 4496) <= temp_inforeg(4511 downto 4504);
					temp_inforeg(4495 downto 4488) <= temp_inforeg(4503 downto 4496);
					temp_inforeg(4487 downto 4480) <= temp_inforeg(4495 downto 4488);
					temp_inforeg(4479 downto 4472) <= temp_inforeg(4487 downto 4480);
					temp_inforeg(4471 downto 4464) <= temp_inforeg(4479 downto 4472);
					temp_inforeg(4463 downto 4456) <= temp_inforeg(4471 downto 4464);
					temp_inforeg(4455 downto 4448) <= temp_inforeg(4463 downto 4456);
					temp_inforeg(4447 downto 4440) <= temp_inforeg(4455 downto 4448);
					temp_inforeg(4439 downto 4432) <= temp_inforeg(4447 downto 4440);
					temp_inforeg(4431 downto 4424) <= temp_inforeg(4439 downto 4432);
					temp_inforeg(4423 downto 4416) <= temp_inforeg(4431 downto 4424);
					temp_inforeg(4415 downto 4408) <= temp_inforeg(4423 downto 4416);
					temp_inforeg(4407 downto 4400) <= temp_inforeg(4415 downto 4408);
					temp_inforeg(4399 downto 4392) <= temp_inforeg(4407 downto 4400);
					temp_inforeg(4391 downto 4384) <= temp_inforeg(4399 downto 4392);
					temp_inforeg(4383 downto 4376) <= temp_inforeg(4391 downto 4384);
					temp_inforeg(4375 downto 4368) <= temp_inforeg(4383 downto 4376);
					temp_inforeg(4367 downto 4360) <= temp_inforeg(4375 downto 4368);
					temp_inforeg(4359 downto 4352) <= temp_inforeg(4367 downto 4360);
					temp_inforeg(4351 downto 4344) <= temp_inforeg(4359 downto 4352);
					temp_inforeg(4343 downto 4336) <= temp_inforeg(4351 downto 4344);
					temp_inforeg(4335 downto 4328) <= temp_inforeg(4343 downto 4336);
					temp_inforeg(4327 downto 4320) <= temp_inforeg(4335 downto 4328);
					temp_inforeg(4319 downto 4312) <= temp_inforeg(4327 downto 4320);
					temp_inforeg(4311 downto 4304) <= temp_inforeg(4319 downto 4312);
					temp_inforeg(4303 downto 4296) <= temp_inforeg(4311 downto 4304);
					temp_inforeg(4295 downto 4288) <= temp_inforeg(4303 downto 4296);
					temp_inforeg(4287 downto 4280) <= temp_inforeg(4295 downto 4288);
					temp_inforeg(4279 downto 4272) <= temp_inforeg(4287 downto 4280);
					temp_inforeg(4271 downto 4264) <= temp_inforeg(4279 downto 4272);
					temp_inforeg(4263 downto 4256) <= temp_inforeg(4271 downto 4264);
					temp_inforeg(4255 downto 4248) <= temp_inforeg(4263 downto 4256);
					temp_inforeg(4247 downto 4240) <= temp_inforeg(4255 downto 4248);
					temp_inforeg(4239 downto 4232) <= temp_inforeg(4247 downto 4240);
					temp_inforeg(4231 downto 4224) <= temp_inforeg(4239 downto 4232);
					temp_inforeg(4223 downto 4216) <= temp_inforeg(4231 downto 4224);
					temp_inforeg(4215 downto 4208) <= temp_inforeg(4223 downto 4216);
					temp_inforeg(4207 downto 4200) <= temp_inforeg(4215 downto 4208);
					temp_inforeg(4199 downto 4192) <= temp_inforeg(4207 downto 4200);
					temp_inforeg(4191 downto 4184) <= temp_inforeg(4199 downto 4192);
					temp_inforeg(4183 downto 4176) <= temp_inforeg(4191 downto 4184);
					temp_inforeg(4175 downto 4168) <= temp_inforeg(4183 downto 4176);
					temp_inforeg(4167 downto 4160) <= temp_inforeg(4175 downto 4168);
					temp_inforeg(4159 downto 4152) <= temp_inforeg(4167 downto 4160);
					temp_inforeg(4151 downto 4144) <= temp_inforeg(4159 downto 4152);
					temp_inforeg(4143 downto 4136) <= temp_inforeg(4151 downto 4144);
					temp_inforeg(4135 downto 4128) <= temp_inforeg(4143 downto 4136);
					temp_inforeg(4127 downto 4120) <= temp_inforeg(4135 downto 4128);
					temp_inforeg(4119 downto 4112) <= temp_inforeg(4127 downto 4120);
					temp_inforeg(4111 downto 4104) <= temp_inforeg(4119 downto 4112);
					temp_inforeg(4103 downto 4096) <= temp_inforeg(4111 downto 4104);
					temp_inforeg(4095 downto 4088) <= temp_inforeg(4103 downto 4096);
					temp_inforeg(4087 downto 4080) <= temp_inforeg(4095 downto 4088);
					temp_inforeg(4079 downto 4072) <= temp_inforeg(4087 downto 4080);
					temp_inforeg(4071 downto 4064) <= temp_inforeg(4079 downto 4072);
					temp_inforeg(4063 downto 4056) <= temp_inforeg(4071 downto 4064);
					temp_inforeg(4055 downto 4048) <= temp_inforeg(4063 downto 4056);
					temp_inforeg(4047 downto 4040) <= temp_inforeg(4055 downto 4048);
					temp_inforeg(4039 downto 4032) <= temp_inforeg(4047 downto 4040);
					temp_inforeg(4031 downto 4024) <= temp_inforeg(4039 downto 4032);
					temp_inforeg(4023 downto 4016) <= temp_inforeg(4031 downto 4024);
					temp_inforeg(4015 downto 4008) <= temp_inforeg(4023 downto 4016);
					temp_inforeg(4007 downto 4000) <= temp_inforeg(4015 downto 4008);
					temp_inforeg(3999 downto 3992) <= temp_inforeg(4007 downto 4000);
					temp_inforeg(3991 downto 3984) <= temp_inforeg(3999 downto 3992);
					temp_inforeg(3983 downto 3976) <= temp_inforeg(3991 downto 3984);
					temp_inforeg(3975 downto 3968) <= temp_inforeg(3983 downto 3976);
					temp_inforeg(3967 downto 3960) <= temp_inforeg(3975 downto 3968);
					temp_inforeg(3959 downto 3952) <= temp_inforeg(3967 downto 3960);
					temp_inforeg(3951 downto 3944) <= temp_inforeg(3959 downto 3952);
					temp_inforeg(3943 downto 3936) <= temp_inforeg(3951 downto 3944);
					temp_inforeg(3935 downto 3928) <= temp_inforeg(3943 downto 3936);
					temp_inforeg(3927 downto 3920) <= temp_inforeg(3935 downto 3928);
					temp_inforeg(3919 downto 3912) <= temp_inforeg(3927 downto 3920);
					temp_inforeg(3911 downto 3904) <= temp_inforeg(3919 downto 3912);
					temp_inforeg(3903 downto 3896) <= temp_inforeg(3911 downto 3904);
					temp_inforeg(3895 downto 3888) <= temp_inforeg(3903 downto 3896);
					temp_inforeg(3887 downto 3880) <= temp_inforeg(3895 downto 3888);
					temp_inforeg(3879 downto 3872) <= temp_inforeg(3887 downto 3880);
					temp_inforeg(3871 downto 3864) <= temp_inforeg(3879 downto 3872);
					temp_inforeg(3863 downto 3856) <= temp_inforeg(3871 downto 3864);
					temp_inforeg(3855 downto 3848) <= temp_inforeg(3863 downto 3856);
					temp_inforeg(3847 downto 3840) <= temp_inforeg(3855 downto 3848);
					temp_inforeg(3839 downto 3832) <= temp_inforeg(3847 downto 3840);
					temp_inforeg(3831 downto 3824) <= temp_inforeg(3839 downto 3832);
					temp_inforeg(3823 downto 3816) <= temp_inforeg(3831 downto 3824);
					temp_inforeg(3815 downto 3808) <= temp_inforeg(3823 downto 3816);
					temp_inforeg(3807 downto 3800) <= temp_inforeg(3815 downto 3808);
					temp_inforeg(3799 downto 3792) <= temp_inforeg(3807 downto 3800);
					temp_inforeg(3791 downto 3784) <= temp_inforeg(3799 downto 3792);
					temp_inforeg(3783 downto 3776) <= temp_inforeg(3791 downto 3784);
					temp_inforeg(3775 downto 3768) <= temp_inforeg(3783 downto 3776);
					temp_inforeg(3767 downto 3760) <= temp_inforeg(3775 downto 3768);
					temp_inforeg(3759 downto 3752) <= temp_inforeg(3767 downto 3760);
					temp_inforeg(3751 downto 3744) <= temp_inforeg(3759 downto 3752);
					temp_inforeg(3743 downto 3736) <= temp_inforeg(3751 downto 3744);
					temp_inforeg(3735 downto 3728) <= temp_inforeg(3743 downto 3736);
					temp_inforeg(3727 downto 3720) <= temp_inforeg(3735 downto 3728);
					temp_inforeg(3719 downto 3712) <= temp_inforeg(3727 downto 3720);
					temp_inforeg(3711 downto 3704) <= temp_inforeg(3719 downto 3712);
					temp_inforeg(3703 downto 3696) <= temp_inforeg(3711 downto 3704);
					temp_inforeg(3695 downto 3688) <= temp_inforeg(3703 downto 3696);
					temp_inforeg(3687 downto 3680) <= temp_inforeg(3695 downto 3688);
					temp_inforeg(3679 downto 3672) <= temp_inforeg(3687 downto 3680);
					temp_inforeg(3671 downto 3664) <= temp_inforeg(3679 downto 3672);
					temp_inforeg(3663 downto 3656) <= temp_inforeg(3671 downto 3664);
					temp_inforeg(3655 downto 3648) <= temp_inforeg(3663 downto 3656);
					temp_inforeg(3647 downto 3640) <= temp_inforeg(3655 downto 3648);
					temp_inforeg(3639 downto 3632) <= temp_inforeg(3647 downto 3640);
					temp_inforeg(3631 downto 3624) <= temp_inforeg(3639 downto 3632);
					temp_inforeg(3623 downto 3616) <= temp_inforeg(3631 downto 3624);
					temp_inforeg(3615 downto 3608) <= temp_inforeg(3623 downto 3616);
					temp_inforeg(3607 downto 3600) <= temp_inforeg(3615 downto 3608);
					temp_inforeg(3599 downto 3592) <= temp_inforeg(3607 downto 3600);
					temp_inforeg(3591 downto 3584) <= temp_inforeg(3599 downto 3592);
					temp_inforeg(3583 downto 3576) <= temp_inforeg(3591 downto 3584);
					temp_inforeg(3575 downto 3568) <= temp_inforeg(3583 downto 3576);
					temp_inforeg(3567 downto 3560) <= temp_inforeg(3575 downto 3568);
					temp_inforeg(3559 downto 3552) <= temp_inforeg(3567 downto 3560);
					temp_inforeg(3551 downto 3544) <= temp_inforeg(3559 downto 3552);
					temp_inforeg(3543 downto 3536) <= temp_inforeg(3551 downto 3544);
					temp_inforeg(3535 downto 3528) <= temp_inforeg(3543 downto 3536);
					temp_inforeg(3527 downto 3520) <= temp_inforeg(3535 downto 3528);
					temp_inforeg(3519 downto 3512) <= temp_inforeg(3527 downto 3520);
					temp_inforeg(3511 downto 3504) <= temp_inforeg(3519 downto 3512);
					temp_inforeg(3503 downto 3496) <= temp_inforeg(3511 downto 3504);
					temp_inforeg(3495 downto 3488) <= temp_inforeg(3503 downto 3496);
					temp_inforeg(3487 downto 3480) <= temp_inforeg(3495 downto 3488);
					temp_inforeg(3479 downto 3472) <= temp_inforeg(3487 downto 3480);
					temp_inforeg(3471 downto 3464) <= temp_inforeg(3479 downto 3472);
					temp_inforeg(3463 downto 3456) <= temp_inforeg(3471 downto 3464);
					temp_inforeg(3455 downto 3448) <= temp_inforeg(3463 downto 3456);
					temp_inforeg(3447 downto 3440) <= temp_inforeg(3455 downto 3448);
					temp_inforeg(3439 downto 3432) <= temp_inforeg(3447 downto 3440);
					temp_inforeg(3431 downto 3424) <= temp_inforeg(3439 downto 3432);
					temp_inforeg(3423 downto 3416) <= temp_inforeg(3431 downto 3424);
					temp_inforeg(3415 downto 3408) <= temp_inforeg(3423 downto 3416);
					temp_inforeg(3407 downto 3400) <= temp_inforeg(3415 downto 3408);
					temp_inforeg(3399 downto 3392) <= temp_inforeg(3407 downto 3400);
					temp_inforeg(3391 downto 3384) <= temp_inforeg(3399 downto 3392);
					temp_inforeg(3383 downto 3376) <= temp_inforeg(3391 downto 3384);
					temp_inforeg(3375 downto 3368) <= temp_inforeg(3383 downto 3376);
					temp_inforeg(3367 downto 3360) <= temp_inforeg(3375 downto 3368);
					temp_inforeg(3359 downto 3352) <= temp_inforeg(3367 downto 3360);
					temp_inforeg(3351 downto 3344) <= temp_inforeg(3359 downto 3352);
					temp_inforeg(3343 downto 3336) <= temp_inforeg(3351 downto 3344);
					temp_inforeg(3335 downto 3328) <= temp_inforeg(3343 downto 3336);
					temp_inforeg(3327 downto 3320) <= temp_inforeg(3335 downto 3328);
					temp_inforeg(3319 downto 3312) <= temp_inforeg(3327 downto 3320);
					temp_inforeg(3311 downto 3304) <= temp_inforeg(3319 downto 3312);
					temp_inforeg(3303 downto 3296) <= temp_inforeg(3311 downto 3304);
					temp_inforeg(3295 downto 3288) <= temp_inforeg(3303 downto 3296);
					temp_inforeg(3287 downto 3280) <= temp_inforeg(3295 downto 3288);
					temp_inforeg(3279 downto 3272) <= temp_inforeg(3287 downto 3280);
					temp_inforeg(3271 downto 3264) <= temp_inforeg(3279 downto 3272);
					temp_inforeg(3263 downto 3256) <= temp_inforeg(3271 downto 3264);
					temp_inforeg(3255 downto 3248) <= temp_inforeg(3263 downto 3256);
					temp_inforeg(3247 downto 3240) <= temp_inforeg(3255 downto 3248);
					temp_inforeg(3239 downto 3232) <= temp_inforeg(3247 downto 3240);
					temp_inforeg(3231 downto 3224) <= temp_inforeg(3239 downto 3232);
					temp_inforeg(3223 downto 3216) <= temp_inforeg(3231 downto 3224);
					temp_inforeg(3215 downto 3208) <= temp_inforeg(3223 downto 3216);
					temp_inforeg(3207 downto 3200) <= temp_inforeg(3215 downto 3208);
					temp_inforeg(3199 downto 3192) <= temp_inforeg(3207 downto 3200);
					temp_inforeg(3191 downto 3184) <= temp_inforeg(3199 downto 3192);
					temp_inforeg(3183 downto 3176) <= temp_inforeg(3191 downto 3184);
					temp_inforeg(3175 downto 3168) <= temp_inforeg(3183 downto 3176);
					temp_inforeg(3167 downto 3160) <= temp_inforeg(3175 downto 3168);
					temp_inforeg(3159 downto 3152) <= temp_inforeg(3167 downto 3160);
					temp_inforeg(3151 downto 3144) <= temp_inforeg(3159 downto 3152);
					temp_inforeg(3143 downto 3136) <= temp_inforeg(3151 downto 3144);
					temp_inforeg(3135 downto 3128) <= temp_inforeg(3143 downto 3136);
					temp_inforeg(3127 downto 3120) <= temp_inforeg(3135 downto 3128);
					temp_inforeg(3119 downto 3112) <= temp_inforeg(3127 downto 3120);
					temp_inforeg(3111 downto 3104) <= temp_inforeg(3119 downto 3112);
					temp_inforeg(3103 downto 3096) <= temp_inforeg(3111 downto 3104);
					temp_inforeg(3095 downto 3088) <= temp_inforeg(3103 downto 3096);
					temp_inforeg(3087 downto 3080) <= temp_inforeg(3095 downto 3088);
					temp_inforeg(3079 downto 3072) <= temp_inforeg(3087 downto 3080);
					temp_inforeg(3071 downto 3064) <= temp_inforeg(3079 downto 3072);
					temp_inforeg(3063 downto 3056) <= temp_inforeg(3071 downto 3064);
					temp_inforeg(3055 downto 3048) <= temp_inforeg(3063 downto 3056);
					temp_inforeg(3047 downto 3040) <= temp_inforeg(3055 downto 3048);
					temp_inforeg(3039 downto 3032) <= temp_inforeg(3047 downto 3040);
					temp_inforeg(3031 downto 3024) <= temp_inforeg(3039 downto 3032);
					temp_inforeg(3023 downto 3016) <= temp_inforeg(3031 downto 3024);
					temp_inforeg(3015 downto 3008) <= temp_inforeg(3023 downto 3016);
					temp_inforeg(3007 downto 3000) <= temp_inforeg(3015 downto 3008);
					temp_inforeg(2999 downto 2992) <= temp_inforeg(3007 downto 3000);
					temp_inforeg(2991 downto 2984) <= temp_inforeg(2999 downto 2992);
					temp_inforeg(2983 downto 2976) <= temp_inforeg(2991 downto 2984);
					temp_inforeg(2975 downto 2968) <= temp_inforeg(2983 downto 2976);
					temp_inforeg(2967 downto 2960) <= temp_inforeg(2975 downto 2968);
					temp_inforeg(2959 downto 2952) <= temp_inforeg(2967 downto 2960);
					temp_inforeg(2951 downto 2944) <= temp_inforeg(2959 downto 2952);
					temp_inforeg(2943 downto 2936) <= temp_inforeg(2951 downto 2944);
					temp_inforeg(2935 downto 2928) <= temp_inforeg(2943 downto 2936);
					temp_inforeg(2927 downto 2920) <= temp_inforeg(2935 downto 2928);
					temp_inforeg(2919 downto 2912) <= temp_inforeg(2927 downto 2920);
					temp_inforeg(2911 downto 2904) <= temp_inforeg(2919 downto 2912);
					temp_inforeg(2903 downto 2896) <= temp_inforeg(2911 downto 2904);
					temp_inforeg(2895 downto 2888) <= temp_inforeg(2903 downto 2896);
					temp_inforeg(2887 downto 2880) <= temp_inforeg(2895 downto 2888);
					temp_inforeg(2879 downto 2872) <= temp_inforeg(2887 downto 2880);
					temp_inforeg(2871 downto 2864) <= temp_inforeg(2879 downto 2872);
					temp_inforeg(2863 downto 2856) <= temp_inforeg(2871 downto 2864);
					temp_inforeg(2855 downto 2848) <= temp_inforeg(2863 downto 2856);
					temp_inforeg(2847 downto 2840) <= temp_inforeg(2855 downto 2848);
					temp_inforeg(2839 downto 2832) <= temp_inforeg(2847 downto 2840);
					temp_inforeg(2831 downto 2824) <= temp_inforeg(2839 downto 2832);
					temp_inforeg(2823 downto 2816) <= temp_inforeg(2831 downto 2824);
					temp_inforeg(2815 downto 2808) <= temp_inforeg(2823 downto 2816);
					temp_inforeg(2807 downto 2800) <= temp_inforeg(2815 downto 2808);
					temp_inforeg(2799 downto 2792) <= temp_inforeg(2807 downto 2800);
					temp_inforeg(2791 downto 2784) <= temp_inforeg(2799 downto 2792);
					temp_inforeg(2783 downto 2776) <= temp_inforeg(2791 downto 2784);
					temp_inforeg(2775 downto 2768) <= temp_inforeg(2783 downto 2776);
					temp_inforeg(2767 downto 2760) <= temp_inforeg(2775 downto 2768);
					temp_inforeg(2759 downto 2752) <= temp_inforeg(2767 downto 2760);
					temp_inforeg(2751 downto 2744) <= temp_inforeg(2759 downto 2752);
					temp_inforeg(2743 downto 2736) <= temp_inforeg(2751 downto 2744);
					temp_inforeg(2735 downto 2728) <= temp_inforeg(2743 downto 2736);
					temp_inforeg(2727 downto 2720) <= temp_inforeg(2735 downto 2728);
					temp_inforeg(2719 downto 2712) <= temp_inforeg(2727 downto 2720);
					temp_inforeg(2711 downto 2704) <= temp_inforeg(2719 downto 2712);
					temp_inforeg(2703 downto 2696) <= temp_inforeg(2711 downto 2704);
					temp_inforeg(2695 downto 2688) <= temp_inforeg(2703 downto 2696);
					temp_inforeg(2687 downto 2680) <= temp_inforeg(2695 downto 2688);
					temp_inforeg(2679 downto 2672) <= temp_inforeg(2687 downto 2680);
					temp_inforeg(2671 downto 2664) <= temp_inforeg(2679 downto 2672);
					temp_inforeg(2663 downto 2656) <= temp_inforeg(2671 downto 2664);
					temp_inforeg(2655 downto 2648) <= temp_inforeg(2663 downto 2656);
					temp_inforeg(2647 downto 2640) <= temp_inforeg(2655 downto 2648);
					temp_inforeg(2639 downto 2632) <= temp_inforeg(2647 downto 2640);
					temp_inforeg(2631 downto 2624) <= temp_inforeg(2639 downto 2632);
					temp_inforeg(2623 downto 2616) <= temp_inforeg(2631 downto 2624);
					temp_inforeg(2615 downto 2608) <= temp_inforeg(2623 downto 2616);
					temp_inforeg(2607 downto 2600) <= temp_inforeg(2615 downto 2608);
					temp_inforeg(2599 downto 2592) <= temp_inforeg(2607 downto 2600);
					temp_inforeg(2591 downto 2584) <= temp_inforeg(2599 downto 2592);
					temp_inforeg(2583 downto 2576) <= temp_inforeg(2591 downto 2584);
					temp_inforeg(2575 downto 2568) <= temp_inforeg(2583 downto 2576);
					temp_inforeg(2567 downto 2560) <= temp_inforeg(2575 downto 2568);
					temp_inforeg(2559 downto 2552) <= temp_inforeg(2567 downto 2560);
					temp_inforeg(2551 downto 2544) <= temp_inforeg(2559 downto 2552);
					temp_inforeg(2543 downto 2536) <= temp_inforeg(2551 downto 2544);
					temp_inforeg(2535 downto 2528) <= temp_inforeg(2543 downto 2536);
					temp_inforeg(2527 downto 2520) <= temp_inforeg(2535 downto 2528);
					temp_inforeg(2519 downto 2512) <= temp_inforeg(2527 downto 2520);
					temp_inforeg(2511 downto 2504) <= temp_inforeg(2519 downto 2512);
					temp_inforeg(2503 downto 2496) <= temp_inforeg(2511 downto 2504);
					temp_inforeg(2495 downto 2488) <= temp_inforeg(2503 downto 2496);
					temp_inforeg(2487 downto 2480) <= temp_inforeg(2495 downto 2488);
					temp_inforeg(2479 downto 2472) <= temp_inforeg(2487 downto 2480);
					temp_inforeg(2471 downto 2464) <= temp_inforeg(2479 downto 2472);
					temp_inforeg(2463 downto 2456) <= temp_inforeg(2471 downto 2464);
					temp_inforeg(2455 downto 2448) <= temp_inforeg(2463 downto 2456);
					temp_inforeg(2447 downto 2440) <= temp_inforeg(2455 downto 2448);
					temp_inforeg(2439 downto 2432) <= temp_inforeg(2447 downto 2440);
					temp_inforeg(2431 downto 2424) <= temp_inforeg(2439 downto 2432);
					temp_inforeg(2423 downto 2416) <= temp_inforeg(2431 downto 2424);
					temp_inforeg(2415 downto 2408) <= temp_inforeg(2423 downto 2416);
					temp_inforeg(2407 downto 2400) <= temp_inforeg(2415 downto 2408);
					temp_inforeg(2399 downto 2392) <= temp_inforeg(2407 downto 2400);
					temp_inforeg(2391 downto 2384) <= temp_inforeg(2399 downto 2392);
					temp_inforeg(2383 downto 2376) <= temp_inforeg(2391 downto 2384);
					temp_inforeg(2375 downto 2368) <= temp_inforeg(2383 downto 2376);
					temp_inforeg(2367 downto 2360) <= temp_inforeg(2375 downto 2368);
					temp_inforeg(2359 downto 2352) <= temp_inforeg(2367 downto 2360);
					temp_inforeg(2351 downto 2344) <= temp_inforeg(2359 downto 2352);
					temp_inforeg(2343 downto 2336) <= temp_inforeg(2351 downto 2344);
					temp_inforeg(2335 downto 2328) <= temp_inforeg(2343 downto 2336);
					temp_inforeg(2327 downto 2320) <= temp_inforeg(2335 downto 2328);
					temp_inforeg(2319 downto 2312) <= temp_inforeg(2327 downto 2320);
					temp_inforeg(2311 downto 2304) <= temp_inforeg(2319 downto 2312);
					temp_inforeg(2303 downto 2296) <= temp_inforeg(2311 downto 2304);
					temp_inforeg(2295 downto 2288) <= temp_inforeg(2303 downto 2296);
					temp_inforeg(2287 downto 2280) <= temp_inforeg(2295 downto 2288);
					temp_inforeg(2279 downto 2272) <= temp_inforeg(2287 downto 2280);
					temp_inforeg(2271 downto 2264) <= temp_inforeg(2279 downto 2272);
					temp_inforeg(2263 downto 2256) <= temp_inforeg(2271 downto 2264);
					temp_inforeg(2255 downto 2248) <= temp_inforeg(2263 downto 2256);
					temp_inforeg(2247 downto 2240) <= temp_inforeg(2255 downto 2248);
					temp_inforeg(2239 downto 2232) <= temp_inforeg(2247 downto 2240);
					temp_inforeg(2231 downto 2224) <= temp_inforeg(2239 downto 2232);
					temp_inforeg(2223 downto 2216) <= temp_inforeg(2231 downto 2224);
					temp_inforeg(2215 downto 2208) <= temp_inforeg(2223 downto 2216);
					temp_inforeg(2207 downto 2200) <= temp_inforeg(2215 downto 2208);
					temp_inforeg(2199 downto 2192) <= temp_inforeg(2207 downto 2200);
					temp_inforeg(2191 downto 2184) <= temp_inforeg(2199 downto 2192);
					temp_inforeg(2183 downto 2176) <= temp_inforeg(2191 downto 2184);
					temp_inforeg(2175 downto 2168) <= temp_inforeg(2183 downto 2176);
					temp_inforeg(2167 downto 2160) <= temp_inforeg(2175 downto 2168);
					temp_inforeg(2159 downto 2152) <= temp_inforeg(2167 downto 2160);
					temp_inforeg(2151 downto 2144) <= temp_inforeg(2159 downto 2152);
					temp_inforeg(2143 downto 2136) <= temp_inforeg(2151 downto 2144);
					temp_inforeg(2135 downto 2128) <= temp_inforeg(2143 downto 2136);
					temp_inforeg(2127 downto 2120) <= temp_inforeg(2135 downto 2128);
					temp_inforeg(2119 downto 2112) <= temp_inforeg(2127 downto 2120);
					temp_inforeg(2111 downto 2104) <= temp_inforeg(2119 downto 2112);
					temp_inforeg(2103 downto 2096) <= temp_inforeg(2111 downto 2104);
					temp_inforeg(2095 downto 2088) <= temp_inforeg(2103 downto 2096);
					temp_inforeg(2087 downto 2080) <= temp_inforeg(2095 downto 2088);
					temp_inforeg(2079 downto 2072) <= temp_inforeg(2087 downto 2080);
					temp_inforeg(2071 downto 2064) <= temp_inforeg(2079 downto 2072);
					temp_inforeg(2063 downto 2056) <= temp_inforeg(2071 downto 2064);
					temp_inforeg(2055 downto 2048) <= temp_inforeg(2063 downto 2056);
					temp_inforeg(2047 downto 2040) <= temp_inforeg(2055 downto 2048);
					temp_inforeg(2039 downto 2032) <= temp_inforeg(2047 downto 2040);
					temp_inforeg(2031 downto 2024) <= temp_inforeg(2039 downto 2032);
					temp_inforeg(2023 downto 2016) <= temp_inforeg(2031 downto 2024);
					temp_inforeg(2015 downto 2008) <= temp_inforeg(2023 downto 2016);
					temp_inforeg(2007 downto 2000) <= temp_inforeg(2015 downto 2008);
					temp_inforeg(1999 downto 1992) <= temp_inforeg(2007 downto 2000);
					temp_inforeg(1991 downto 1984) <= temp_inforeg(1999 downto 1992);
					temp_inforeg(1983 downto 1976) <= temp_inforeg(1991 downto 1984);
					temp_inforeg(1975 downto 1968) <= temp_inforeg(1983 downto 1976);
					temp_inforeg(1967 downto 1960) <= temp_inforeg(1975 downto 1968);
					temp_inforeg(1959 downto 1952) <= temp_inforeg(1967 downto 1960);
					temp_inforeg(1951 downto 1944) <= temp_inforeg(1959 downto 1952);
					temp_inforeg(1943 downto 1936) <= temp_inforeg(1951 downto 1944);
					temp_inforeg(1935 downto 1928) <= temp_inforeg(1943 downto 1936);
					temp_inforeg(1927 downto 1920) <= temp_inforeg(1935 downto 1928);
					temp_inforeg(1919 downto 1912) <= temp_inforeg(1927 downto 1920);
					temp_inforeg(1911 downto 1904) <= temp_inforeg(1919 downto 1912);
					temp_inforeg(1903 downto 1896) <= temp_inforeg(1911 downto 1904);
					temp_inforeg(1895 downto 1888) <= temp_inforeg(1903 downto 1896);
					temp_inforeg(1887 downto 1880) <= temp_inforeg(1895 downto 1888);
					temp_inforeg(1879 downto 1872) <= temp_inforeg(1887 downto 1880);
					temp_inforeg(1871 downto 1864) <= temp_inforeg(1879 downto 1872);
					temp_inforeg(1863 downto 1856) <= temp_inforeg(1871 downto 1864);
					temp_inforeg(1855 downto 1848) <= temp_inforeg(1863 downto 1856);
					temp_inforeg(1847 downto 1840) <= temp_inforeg(1855 downto 1848);
					temp_inforeg(1839 downto 1832) <= temp_inforeg(1847 downto 1840);
					temp_inforeg(1831 downto 1824) <= temp_inforeg(1839 downto 1832);
					temp_inforeg(1823 downto 1816) <= temp_inforeg(1831 downto 1824);
					temp_inforeg(1815 downto 1808) <= temp_inforeg(1823 downto 1816);
					temp_inforeg(1807 downto 1800) <= temp_inforeg(1815 downto 1808);
					temp_inforeg(1799 downto 1792) <= temp_inforeg(1807 downto 1800);
					temp_inforeg(1791 downto 1784) <= temp_inforeg(1799 downto 1792);
					temp_inforeg(1783 downto 1776) <= temp_inforeg(1791 downto 1784);
					temp_inforeg(1775 downto 1768) <= temp_inforeg(1783 downto 1776);
					temp_inforeg(1767 downto 1760) <= temp_inforeg(1775 downto 1768);
					temp_inforeg(1759 downto 1752) <= temp_inforeg(1767 downto 1760);
					temp_inforeg(1751 downto 1744) <= temp_inforeg(1759 downto 1752);
					temp_inforeg(1743 downto 1736) <= temp_inforeg(1751 downto 1744);
					temp_inforeg(1735 downto 1728) <= temp_inforeg(1743 downto 1736);
					temp_inforeg(1727 downto 1720) <= temp_inforeg(1735 downto 1728);
					temp_inforeg(1719 downto 1712) <= temp_inforeg(1727 downto 1720);
					temp_inforeg(1711 downto 1704) <= temp_inforeg(1719 downto 1712);
					temp_inforeg(1703 downto 1696) <= temp_inforeg(1711 downto 1704);
					temp_inforeg(1695 downto 1688) <= temp_inforeg(1703 downto 1696);
					temp_inforeg(1687 downto 1680) <= temp_inforeg(1695 downto 1688);
					temp_inforeg(1679 downto 1672) <= temp_inforeg(1687 downto 1680);
					temp_inforeg(1671 downto 1664) <= temp_inforeg(1679 downto 1672);
					temp_inforeg(1663 downto 1656) <= temp_inforeg(1671 downto 1664);
					temp_inforeg(1655 downto 1648) <= temp_inforeg(1663 downto 1656);
					temp_inforeg(1647 downto 1640) <= temp_inforeg(1655 downto 1648);
					temp_inforeg(1639 downto 1632) <= temp_inforeg(1647 downto 1640);
					temp_inforeg(1631 downto 1624) <= temp_inforeg(1639 downto 1632);
					temp_inforeg(1623 downto 1616) <= temp_inforeg(1631 downto 1624);
					temp_inforeg(1615 downto 1608) <= temp_inforeg(1623 downto 1616);
					temp_inforeg(1607 downto 1600) <= temp_inforeg(1615 downto 1608);
					temp_inforeg(1599 downto 1592) <= temp_inforeg(1607 downto 1600);
					temp_inforeg(1591 downto 1584) <= temp_inforeg(1599 downto 1592);
					temp_inforeg(1583 downto 1576) <= temp_inforeg(1591 downto 1584);
					temp_inforeg(1575 downto 1568) <= temp_inforeg(1583 downto 1576);
					temp_inforeg(1567 downto 1560) <= temp_inforeg(1575 downto 1568);
					temp_inforeg(1559 downto 1552) <= temp_inforeg(1567 downto 1560);
					temp_inforeg(1551 downto 1544) <= temp_inforeg(1559 downto 1552);
					temp_inforeg(1543 downto 1536) <= temp_inforeg(1551 downto 1544);
					temp_inforeg(1535 downto 1528) <= temp_inforeg(1543 downto 1536);
					temp_inforeg(1527 downto 1520) <= temp_inforeg(1535 downto 1528);
					temp_inforeg(1519 downto 1512) <= temp_inforeg(1527 downto 1520);
					temp_inforeg(1511 downto 1504) <= temp_inforeg(1519 downto 1512);
					temp_inforeg(1503 downto 1496) <= temp_inforeg(1511 downto 1504);
					temp_inforeg(1495 downto 1488) <= temp_inforeg(1503 downto 1496);
					temp_inforeg(1487 downto 1480) <= temp_inforeg(1495 downto 1488);
					temp_inforeg(1479 downto 1472) <= temp_inforeg(1487 downto 1480);
					temp_inforeg(1471 downto 1464) <= temp_inforeg(1479 downto 1472);
					temp_inforeg(1463 downto 1456) <= temp_inforeg(1471 downto 1464);
					temp_inforeg(1455 downto 1448) <= temp_inforeg(1463 downto 1456);
					temp_inforeg(1447 downto 1440) <= temp_inforeg(1455 downto 1448);
					temp_inforeg(1439 downto 1432) <= temp_inforeg(1447 downto 1440);
					temp_inforeg(1431 downto 1424) <= temp_inforeg(1439 downto 1432);
					temp_inforeg(1423 downto 1416) <= temp_inforeg(1431 downto 1424);
					temp_inforeg(1415 downto 1408) <= temp_inforeg(1423 downto 1416);
					temp_inforeg(1407 downto 1400) <= temp_inforeg(1415 downto 1408);
					temp_inforeg(1399 downto 1392) <= temp_inforeg(1407 downto 1400);
					temp_inforeg(1391 downto 1384) <= temp_inforeg(1399 downto 1392);
					temp_inforeg(1383 downto 1376) <= temp_inforeg(1391 downto 1384);
					temp_inforeg(1375 downto 1368) <= temp_inforeg(1383 downto 1376);
					temp_inforeg(1367 downto 1360) <= temp_inforeg(1375 downto 1368);
					temp_inforeg(1359 downto 1352) <= temp_inforeg(1367 downto 1360);
					temp_inforeg(1351 downto 1344) <= temp_inforeg(1359 downto 1352);
					temp_inforeg(1343 downto 1336) <= temp_inforeg(1351 downto 1344);
					temp_inforeg(1335 downto 1328) <= temp_inforeg(1343 downto 1336);
					temp_inforeg(1327 downto 1320) <= temp_inforeg(1335 downto 1328);
					temp_inforeg(1319 downto 1312) <= temp_inforeg(1327 downto 1320);
					temp_inforeg(1311 downto 1304) <= temp_inforeg(1319 downto 1312);
					temp_inforeg(1303 downto 1296) <= temp_inforeg(1311 downto 1304);
					temp_inforeg(1295 downto 1288) <= temp_inforeg(1303 downto 1296);
					temp_inforeg(1287 downto 1280) <= temp_inforeg(1295 downto 1288);
					temp_inforeg(1279 downto 1272) <= temp_inforeg(1287 downto 1280);
					temp_inforeg(1271 downto 1264) <= temp_inforeg(1279 downto 1272);
					temp_inforeg(1263 downto 1256) <= temp_inforeg(1271 downto 1264);
					temp_inforeg(1255 downto 1248) <= temp_inforeg(1263 downto 1256);
					temp_inforeg(1247 downto 1240) <= temp_inforeg(1255 downto 1248);
					temp_inforeg(1239 downto 1232) <= temp_inforeg(1247 downto 1240);
					temp_inforeg(1231 downto 1224) <= temp_inforeg(1239 downto 1232);
					temp_inforeg(1223 downto 1216) <= temp_inforeg(1231 downto 1224);
					temp_inforeg(1215 downto 1208) <= temp_inforeg(1223 downto 1216);
					temp_inforeg(1207 downto 1200) <= temp_inforeg(1215 downto 1208);
					temp_inforeg(1199 downto 1192) <= temp_inforeg(1207 downto 1200);
					temp_inforeg(1191 downto 1184) <= temp_inforeg(1199 downto 1192);
					temp_inforeg(1183 downto 1176) <= temp_inforeg(1191 downto 1184);
					temp_inforeg(1175 downto 1168) <= temp_inforeg(1183 downto 1176);
					temp_inforeg(1167 downto 1160) <= temp_inforeg(1175 downto 1168);
					temp_inforeg(1159 downto 1152) <= temp_inforeg(1167 downto 1160);
					temp_inforeg(1151 downto 1144) <= temp_inforeg(1159 downto 1152);
					temp_inforeg(1143 downto 1136) <= temp_inforeg(1151 downto 1144);
					temp_inforeg(1135 downto 1128) <= temp_inforeg(1143 downto 1136);
					temp_inforeg(1127 downto 1120) <= temp_inforeg(1135 downto 1128);
					temp_inforeg(1119 downto 1112) <= temp_inforeg(1127 downto 1120);
					temp_inforeg(1111 downto 1104) <= temp_inforeg(1119 downto 1112);
					temp_inforeg(1103 downto 1096) <= temp_inforeg(1111 downto 1104);
					temp_inforeg(1095 downto 1088) <= temp_inforeg(1103 downto 1096);
					temp_inforeg(1087 downto 1080) <= temp_inforeg(1095 downto 1088);
					temp_inforeg(1079 downto 1072) <= temp_inforeg(1087 downto 1080);
					temp_inforeg(1071 downto 1064) <= temp_inforeg(1079 downto 1072);
					temp_inforeg(1063 downto 1056) <= temp_inforeg(1071 downto 1064);
					temp_inforeg(1055 downto 1048) <= temp_inforeg(1063 downto 1056);
					temp_inforeg(1047 downto 1040) <= temp_inforeg(1055 downto 1048);
					temp_inforeg(1039 downto 1032) <= temp_inforeg(1047 downto 1040);
					temp_inforeg(1031 downto 1024) <= temp_inforeg(1039 downto 1032);
					temp_inforeg(1023 downto 1016) <= temp_inforeg(1031 downto 1024);
					temp_inforeg(1015 downto 1008) <= temp_inforeg(1023 downto 1016);
					temp_inforeg(1007 downto 1000) <= temp_inforeg(1015 downto 1008);
					temp_inforeg(999 downto 992) <= temp_inforeg(1007 downto 1000);
					temp_inforeg(991 downto 984) <= temp_inforeg(999 downto 992);
					temp_inforeg(983 downto 976) <= temp_inforeg(991 downto 984);
					temp_inforeg(975 downto 968) <= temp_inforeg(983 downto 976);
					temp_inforeg(967 downto 960) <= temp_inforeg(975 downto 968);
					temp_inforeg(959 downto 952) <= temp_inforeg(967 downto 960);
					temp_inforeg(951 downto 944) <= temp_inforeg(959 downto 952);
					temp_inforeg(943 downto 936) <= temp_inforeg(951 downto 944);
					temp_inforeg(935 downto 928) <= temp_inforeg(943 downto 936);
					temp_inforeg(927 downto 920) <= temp_inforeg(935 downto 928);
					temp_inforeg(919 downto 912) <= temp_inforeg(927 downto 920);
					temp_inforeg(911 downto 904) <= temp_inforeg(919 downto 912);
					temp_inforeg(903 downto 896) <= temp_inforeg(911 downto 904);
					temp_inforeg(895 downto 888) <= temp_inforeg(903 downto 896);
					temp_inforeg(887 downto 880) <= temp_inforeg(895 downto 888);
					temp_inforeg(879 downto 872) <= temp_inforeg(887 downto 880);
					temp_inforeg(871 downto 864) <= temp_inforeg(879 downto 872);
					temp_inforeg(863 downto 856) <= temp_inforeg(871 downto 864);
					temp_inforeg(855 downto 848) <= temp_inforeg(863 downto 856);
					temp_inforeg(847 downto 840) <= temp_inforeg(855 downto 848);
					temp_inforeg(839 downto 832) <= temp_inforeg(847 downto 840);
					temp_inforeg(831 downto 824) <= temp_inforeg(839 downto 832);
					temp_inforeg(823 downto 816) <= temp_inforeg(831 downto 824);
					temp_inforeg(815 downto 808) <= temp_inforeg(823 downto 816);
					temp_inforeg(807 downto 800) <= temp_inforeg(815 downto 808);
					temp_inforeg(799 downto 792) <= temp_inforeg(807 downto 800);
					temp_inforeg(791 downto 784) <= temp_inforeg(799 downto 792);
					temp_inforeg(783 downto 776) <= temp_inforeg(791 downto 784);
					temp_inforeg(775 downto 768) <= temp_inforeg(783 downto 776);
					temp_inforeg(767 downto 760) <= temp_inforeg(775 downto 768);
					temp_inforeg(759 downto 752) <= temp_inforeg(767 downto 760);
					temp_inforeg(751 downto 744) <= temp_inforeg(759 downto 752);
					temp_inforeg(743 downto 736) <= temp_inforeg(751 downto 744);
					temp_inforeg(735 downto 728) <= temp_inforeg(743 downto 736);
					temp_inforeg(727 downto 720) <= temp_inforeg(735 downto 728);
					temp_inforeg(719 downto 712) <= temp_inforeg(727 downto 720);
					temp_inforeg(711 downto 704) <= temp_inforeg(719 downto 712);
					temp_inforeg(703 downto 696) <= temp_inforeg(711 downto 704);
					temp_inforeg(695 downto 688) <= temp_inforeg(703 downto 696);
					temp_inforeg(687 downto 680) <= temp_inforeg(695 downto 688);
					temp_inforeg(679 downto 672) <= temp_inforeg(687 downto 680);
					temp_inforeg(671 downto 664) <= temp_inforeg(679 downto 672);
					temp_inforeg(663 downto 656) <= temp_inforeg(671 downto 664);
					temp_inforeg(655 downto 648) <= temp_inforeg(663 downto 656);
					temp_inforeg(647 downto 640) <= temp_inforeg(655 downto 648);
					temp_inforeg(639 downto 632) <= temp_inforeg(647 downto 640);
					temp_inforeg(631 downto 624) <= temp_inforeg(639 downto 632);
					temp_inforeg(623 downto 616) <= temp_inforeg(631 downto 624);
					temp_inforeg(615 downto 608) <= temp_inforeg(623 downto 616);
					temp_inforeg(607 downto 600) <= temp_inforeg(615 downto 608);
					temp_inforeg(599 downto 592) <= temp_inforeg(607 downto 600);
					temp_inforeg(591 downto 584) <= temp_inforeg(599 downto 592);
					temp_inforeg(583 downto 576) <= temp_inforeg(591 downto 584);
					temp_inforeg(575 downto 568) <= temp_inforeg(583 downto 576);
					temp_inforeg(567 downto 560) <= temp_inforeg(575 downto 568);
					temp_inforeg(559 downto 552) <= temp_inforeg(567 downto 560);
					temp_inforeg(551 downto 544) <= temp_inforeg(559 downto 552);
					temp_inforeg(543 downto 536) <= temp_inforeg(551 downto 544);
					temp_inforeg(535 downto 528) <= temp_inforeg(543 downto 536);
					temp_inforeg(527 downto 520) <= temp_inforeg(535 downto 528);
					temp_inforeg(519 downto 512) <= temp_inforeg(527 downto 520);
					temp_inforeg(511 downto 504) <= temp_inforeg(519 downto 512);
					temp_inforeg(503 downto 496) <= temp_inforeg(511 downto 504);
					temp_inforeg(495 downto 488) <= temp_inforeg(503 downto 496);
					temp_inforeg(487 downto 480) <= temp_inforeg(495 downto 488);
					temp_inforeg(479 downto 472) <= temp_inforeg(487 downto 480);
					temp_inforeg(471 downto 464) <= temp_inforeg(479 downto 472);
					temp_inforeg(463 downto 456) <= temp_inforeg(471 downto 464);
					temp_inforeg(455 downto 448) <= temp_inforeg(463 downto 456);
					temp_inforeg(447 downto 440) <= temp_inforeg(455 downto 448);
					temp_inforeg(439 downto 432) <= temp_inforeg(447 downto 440);
					temp_inforeg(431 downto 424) <= temp_inforeg(439 downto 432);
					temp_inforeg(423 downto 416) <= temp_inforeg(431 downto 424);
					temp_inforeg(415 downto 408) <= temp_inforeg(423 downto 416);
					temp_inforeg(407 downto 400) <= temp_inforeg(415 downto 408);
					temp_inforeg(399 downto 392) <= temp_inforeg(407 downto 400);
					temp_inforeg(391 downto 384) <= temp_inforeg(399 downto 392);
					temp_inforeg(383 downto 376) <= temp_inforeg(391 downto 384);
					temp_inforeg(375 downto 368) <= temp_inforeg(383 downto 376);
					temp_inforeg(367 downto 360) <= temp_inforeg(375 downto 368);
					temp_inforeg(359 downto 352) <= temp_inforeg(367 downto 360);
					temp_inforeg(351 downto 344) <= temp_inforeg(359 downto 352);
					temp_inforeg(343 downto 336) <= temp_inforeg(351 downto 344);
					temp_inforeg(335 downto 328) <= temp_inforeg(343 downto 336);
					temp_inforeg(327 downto 320) <= temp_inforeg(335 downto 328);
					temp_inforeg(319 downto 312) <= temp_inforeg(327 downto 320);
					temp_inforeg(311 downto 304) <= temp_inforeg(319 downto 312);
					temp_inforeg(303 downto 296) <= temp_inforeg(311 downto 304);
					temp_inforeg(295 downto 288) <= temp_inforeg(303 downto 296);
					temp_inforeg(287 downto 280) <= temp_inforeg(295 downto 288);
					temp_inforeg(279 downto 272) <= temp_inforeg(287 downto 280);
					temp_inforeg(271 downto 264) <= temp_inforeg(279 downto 272);
					temp_inforeg(263 downto 256) <= temp_inforeg(271 downto 264);
					temp_inforeg(255 downto 248) <= temp_inforeg(263 downto 256);
					temp_inforeg(247 downto 240) <= temp_inforeg(255 downto 248);
					temp_inforeg(239 downto 232) <= temp_inforeg(247 downto 240);
					temp_inforeg(231 downto 224) <= temp_inforeg(239 downto 232);
					temp_inforeg(223 downto 216) <= temp_inforeg(231 downto 224);
					temp_inforeg(215 downto 208) <= temp_inforeg(223 downto 216);
					temp_inforeg(207 downto 200) <= temp_inforeg(215 downto 208);
					temp_inforeg(199 downto 192) <= temp_inforeg(207 downto 200);
					temp_inforeg(191 downto 184) <= temp_inforeg(199 downto 192);
					temp_inforeg(183 downto 176) <= temp_inforeg(191 downto 184);
					temp_inforeg(175 downto 168) <= temp_inforeg(183 downto 176);
					temp_inforeg(167 downto 160) <= temp_inforeg(175 downto 168);
					temp_inforeg(159 downto 152) <= temp_inforeg(167 downto 160);
					temp_inforeg(151 downto 144) <= temp_inforeg(159 downto 152);
					temp_inforeg(143 downto 136) <= temp_inforeg(151 downto 144);
					temp_inforeg(135 downto 128) <= temp_inforeg(143 downto 136);
					temp_inforeg(127 downto 120) <= temp_inforeg(135 downto 128);
					temp_inforeg(119 downto 112) <= temp_inforeg(127 downto 120);
					temp_inforeg(111 downto 104) <= temp_inforeg(119 downto 112);
					temp_inforeg(103 downto 96) <= temp_inforeg(111 downto 104);
					temp_inforeg(95 downto 88) <= temp_inforeg(103 downto 96);
					temp_inforeg(87 downto 80) <= temp_inforeg(95 downto 88);
					temp_inforeg(79 downto 72) <= temp_inforeg(87 downto 80);
					temp_inforeg(71 downto 64) <= temp_inforeg(79 downto 72);
					temp_inforeg(63 downto 56) <= temp_inforeg(71 downto 64);
					temp_inforeg(55 downto 48) <= temp_inforeg(63 downto 56);
					temp_inforeg(47 downto 40) <= temp_inforeg(55 downto 48);
					temp_inforeg(39 downto 32) <= temp_inforeg(47 downto 40);
					temp_inforeg(31 downto 24) <= temp_inforeg(39 downto 32);
					temp_inforeg(23 downto 16) <= temp_inforeg(31 downto 24);
					temp_inforeg(15 downto 8) <= temp_inforeg(23 downto 16);
					temp_inforeg(7 downto 0) <= temp_inforeg(15 downto 8);
				end if;
			end if;
		end process;
	end rtl;
