lvds_tx_DA_inst : lvds_tx_DA PORT MAP (
		tx_in	 => tx_in_sig,
		tx_inclock	 => tx_inclock_sig,
		tx_out	 => tx_out_sig
	);
